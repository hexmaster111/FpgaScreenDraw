/* verilator lint_off UNDRIVEN */
/* verilator lint_off UNUSEDSIGNAL */
/* verilator lint_off UNUSEDPARAM */
module videomem2 (
    input  wire [9:0] vm_px, vm_py, // px being scanned right now
    input  wire [7:0] vm_ch_in,
    input  wire       vm_ch_write_enable, write_clk,
    output wire [5:0] vm_r, vm_g, vm_b, // output rgb colors
    output wire [7:0] debug_curr_ch_out
);

parameter DISP_WIDTH_PX  = 640;
parameter DISP_HEIGHT_PX = 480;
parameter CH_WIDTH = 4;
parameter CH_HEIGHT = 8;
parameter CH_WIDTH_SCREEN = DISP_WIDTH_PX / CH_WIDTH;
parameter CH_HEIGHT_SCREEN = DISP_HEIGHT_PX / CH_HEIGHT;
parameter CH_SCREENSIZE = CH_WIDTH_SCREEN * CH_HEIGHT_SCREEN;

  // 640 x 480 px screen size
  // 160 x  60 chars on screen 
  //   4 x   8 px char size
  //      9600 chars in video memory
reg [7:0] vmem [CH_SCREENSIZE-1:0]; // 9600x  8 bit values


wire  [7:0] char_out;
wire [31:0] char_gfx;
fontrom fr(char_out, char_gfx);


assign char_out = vmem [(vm_py / CH_HEIGHT) * CH_WIDTH_SCREEN + (vm_px / CH_WIDTH)];
// assign char_out = 8'd87;
assign debug_curr_ch_out = char_out;
//abcdefghijklmnopqrstuvwxyz

/*
char_x_px = vm_px / CH_WIDTH;
char_y_px = vm_py / CH_HEIGHT;
bit = char_y_px * CH_WIDTH + char_x_px;
r g b = bit ? 1 : 0

                int bit = (gfx >> (y * 4 + x)) & 1; 
*/
assign vm_r = char_gfx[((vm_py % CH_HEIGHT) * CH_WIDTH) + (vm_px % CH_WIDTH)] ? 6'b111111 : 6'b000000;
assign vm_g = char_gfx[((vm_py % CH_HEIGHT) * CH_WIDTH) + (vm_px % CH_WIDTH)] ? 6'b111111 : 6'b000000;
assign vm_b = char_gfx[((vm_py % CH_HEIGHT) * CH_WIDTH) + (vm_px % CH_WIDTH)] ? 6'b111111 : 6'b000000;

always @(posedge write_clk) begin
    if(vm_ch_write_enable == 1'b1) begin // write
        // todo : write into vmem
    end
end

integer i;
initial begin
    
    // lol quartus just wouldnt let it itterate more then 5000 times
    for (i = 0; i < CH_SCREENSIZE/2; i = i + 1) begin
        vmem[i] = 8'd32; // ASCII for space ' '
    end

    for (i = CH_SCREENSIZE/2; i < CH_SCREENSIZE; i = i + 1) begin
        vmem[i] = 8'd32; // ASCII for space ' '
    end

    for (i = 0; i < 255; i = i + 1) begin
        vmem[i] = i; // ASCII for space ' '
    end

    
vmem[258] = 8'd116;
vmem[259] = 8'd105;
vmem[260] = 8'd97;
vmem[261] = 8'd109;
vmem[262] = 8'd32;
vmem[263] = 8'd102;
vmem[264] = 8'd101;
vmem[265] = 8'd114;
vmem[266] = 8'd109;
vmem[267] = 8'd101;
vmem[268] = 8'd110;
vmem[269] = 8'd116;
vmem[270] = 8'd117;
vmem[271] = 8'd109;
vmem[272] = 8'd32;
vmem[273] = 8'd110;
vmem[274] = 8'd101;
vmem[275] = 8'd99;
vmem[276] = 8'd32;
vmem[277] = 8'd112;
vmem[278] = 8'd117;
vmem[279] = 8'd114;
vmem[280] = 8'd117;
vmem[281] = 8'd115;
vmem[282] = 8'd32;
vmem[283] = 8'd101;
vmem[284] = 8'd116;
vmem[285] = 8'd32;
vmem[286] = 8'd112;
vmem[287] = 8'd117;
vmem[288] = 8'd108;
vmem[289] = 8'd118;
vmem[290] = 8'd105;
vmem[291] = 8'd110;
vmem[292] = 8'd97;
vmem[293] = 8'd114;
vmem[294] = 8'd46;
vmem[295] = 8'd32;
vmem[296] = 8'd78;
vmem[297] = 8'd97;
vmem[298] = 8'd109;
vmem[299] = 8'd32;
vmem[300] = 8'd115;
vmem[301] = 8'd111;
vmem[302] = 8'd100;
vmem[303] = 8'd97;
vmem[304] = 8'd108;
vmem[305] = 8'd101;
vmem[306] = 8'd115;
vmem[307] = 8'd32;
vmem[308] = 8'd116;
vmem[309] = 8'd101;
vmem[310] = 8'd109;
vmem[311] = 8'd112;
vmem[312] = 8'd111;
vmem[313] = 8'd114;
vmem[314] = 8'd32;
vmem[315] = 8'd109;
vmem[316] = 8'd105;
vmem[317] = 8'd32;
vmem[318] = 8'd101;
vmem[319] = 8'd103;
vmem[320] = 8'd101;
vmem[321] = 8'd116;
vmem[322] = 8'd32;
vmem[323] = 8'd109;
vmem[324] = 8'd97;
vmem[325] = 8'd120;
vmem[326] = 8'd105;
vmem[327] = 8'd109;
vmem[328] = 8'd117;
vmem[329] = 8'd115;
vmem[330] = 8'd46;
vmem[331] = 8'd32;
vmem[332] = 8'd67;
vmem[333] = 8'd114;
vmem[334] = 8'd97;
vmem[335] = 8'd115;
vmem[336] = 8'd32;
vmem[337] = 8'd98;
vmem[338] = 8'd108;
vmem[339] = 8'd97;
vmem[340] = 8'd110;
vmem[341] = 8'd100;
vmem[342] = 8'd105;
vmem[343] = 8'd116;
vmem[344] = 8'd32;
vmem[345] = 8'd97;
vmem[346] = 8'd99;
vmem[347] = 8'd32;
vmem[348] = 8'd109;
vmem[349] = 8'd97;
vmem[350] = 8'd103;
vmem[351] = 8'd110;
vmem[352] = 8'd97;
vmem[353] = 8'd32;
vmem[354] = 8'd115;
vmem[355] = 8'd101;
vmem[356] = 8'd100;
vmem[357] = 8'd32;
vmem[358] = 8'd112;
vmem[359] = 8'd111;
vmem[360] = 8'd115;
vmem[361] = 8'd117;
vmem[362] = 8'd101;
vmem[363] = 8'd114;
vmem[364] = 8'd101;
vmem[365] = 8'd46;
vmem[366] = 8'd32;
vmem[367] = 8'd77;
vmem[368] = 8'd97;
vmem[369] = 8'd101;
vmem[370] = 8'd99;
vmem[371] = 8'd101;
vmem[372] = 8'd110;
vmem[373] = 8'd97;
vmem[374] = 8'd115;
vmem[375] = 8'd32;
vmem[376] = 8'd100;
vmem[377] = 8'd105;
vmem[378] = 8'd103;
vmem[379] = 8'd110;
vmem[380] = 8'd105;
vmem[381] = 8'd115;
vmem[382] = 8'd115;
vmem[383] = 8'd105;
vmem[384] = 8'd109;
vmem[385] = 8'd44;
vmem[386] = 8'd32;
vmem[387] = 8'd109;
vmem[388] = 8'd97;
vmem[389] = 8'd115;
vmem[390] = 8'd115;
vmem[391] = 8'd97;
vmem[392] = 8'd32;
vmem[393] = 8'd113;
vmem[394] = 8'd117;
vmem[395] = 8'd105;
vmem[396] = 8'd115;
vmem[397] = 8'd32;
vmem[398] = 8'd116;
vmem[399] = 8'd101;
vmem[400] = 8'd109;
vmem[401] = 8'd112;
vmem[402] = 8'd111;
vmem[403] = 8'd114;
vmem[404] = 8'd32;
vmem[405] = 8'd105;
vmem[406] = 8'd97;
vmem[407] = 8'd99;
vmem[408] = 8'd117;
vmem[409] = 8'd108;
vmem[410] = 8'd105;
vmem[411] = 8'd115;
vmem[412] = 8'd44;
vmem[413] = 8'd32;
vmem[414] = 8'd114;
vmem[415] = 8'd105;
vmem[416] = 8'd115;
vmem[417] = 8'd117;
vmem[418] = 8'd115;
vmem[419] = 8'd32;
vmem[420] = 8'd97;
vmem[421] = 8'd114;
vmem[422] = 8'd99;
vmem[423] = 8'd117;
vmem[424] = 8'd32;
vmem[425] = 8'd98;
vmem[426] = 8'd108;
vmem[427] = 8'd97;
vmem[428] = 8'd110;
vmem[429] = 8'd100;
vmem[430] = 8'd105;
vmem[431] = 8'd116;
vmem[432] = 8'd32;
vmem[433] = 8'd101;
vmem[434] = 8'd108;
vmem[435] = 8'd105;
vmem[436] = 8'd116;
vmem[437] = 8'd44;
vmem[438] = 8'd32;
vmem[439] = 8'd110;
vmem[440] = 8'd111;
vmem[441] = 8'd110;
vmem[442] = 8'd32;
vmem[443] = 8'd109;
vmem[444] = 8'd111;
vmem[445] = 8'd108;
vmem[446] = 8'd108;
vmem[447] = 8'd105;
vmem[448] = 8'd115;
vmem[449] = 8'd32;
vmem[450] = 8'd110;
vmem[451] = 8'd117;
vmem[452] = 8'd110;
vmem[453] = 8'd99;
vmem[454] = 8'd32;
vmem[455] = 8'd116;
vmem[456] = 8'd101;
vmem[457] = 8'd108;
vmem[458] = 8'd108;
vmem[459] = 8'd117;
vmem[460] = 8'd115;
vmem[461] = 8'd32;
vmem[462] = 8'd100;
vmem[463] = 8'd97;
vmem[464] = 8'd112;
vmem[465] = 8'd105;
vmem[466] = 8'd98;
vmem[467] = 8'd117;
vmem[468] = 8'd115;
vmem[469] = 8'd32;
vmem[470] = 8'd109;
vmem[471] = 8'd105;
vmem[472] = 8'd46;
vmem[473] = 8'd32;
vmem[474] = 8'd67;
vmem[475] = 8'd117;
vmem[476] = 8'd114;
vmem[477] = 8'd97;
vmem[478] = 8'd98;
vmem[479] = 8'd105;
vmem[480] = 8'd116;
vmem[481] = 8'd117;
vmem[482] = 8'd114;
vmem[483] = 8'd32;
vmem[484] = 8'd112;
vmem[485] = 8'd117;
vmem[486] = 8'd108;
vmem[487] = 8'd118;
vmem[488] = 8'd105;
vmem[489] = 8'd110;
vmem[490] = 8'd97;
vmem[491] = 8'd114;
vmem[492] = 8'd32;
vmem[493] = 8'd100;
vmem[494] = 8'd117;
vmem[495] = 8'd105;
vmem[496] = 8'd32;
vmem[497] = 8'd115;
vmem[498] = 8'd101;
vmem[499] = 8'd100;
vmem[500] = 8'd32;
vmem[501] = 8'd102;
vmem[502] = 8'd97;
vmem[503] = 8'd99;
vmem[504] = 8'd105;
vmem[505] = 8'd108;
vmem[506] = 8'd105;
vmem[507] = 8'd115;
vmem[508] = 8'd105;
vmem[509] = 8'd115;
vmem[510] = 8'd32;
vmem[511] = 8'd118;
vmem[512] = 8'd101;
vmem[513] = 8'd104;
vmem[514] = 8'd105;
vmem[515] = 8'd99;
vmem[516] = 8'd117;
vmem[517] = 8'd108;
vmem[518] = 8'd97;
vmem[519] = 8'd46;
vmem[520] = 8'd32;
vmem[521] = 8'd67;
vmem[522] = 8'd114;
vmem[523] = 8'd97;
vmem[524] = 8'd115;
vmem[525] = 8'd32;
vmem[526] = 8'd117;
vmem[527] = 8'd116;
vmem[528] = 8'd32;
vmem[529] = 8'd114;
vmem[530] = 8'd105;
vmem[531] = 8'd115;
vmem[532] = 8'd117;
vmem[533] = 8'd115;
vmem[534] = 8'd32;
vmem[535] = 8'd110;
vmem[536] = 8'd101;
vmem[537] = 8'd113;
vmem[538] = 8'd117;
vmem[539] = 8'd101;
vmem[540] = 8'd46;
vmem[541] = 8'd32;
vmem[542] = 8'd67;
vmem[543] = 8'd117;
vmem[544] = 8'd114;
vmem[545] = 8'd97;
vmem[546] = 8'd98;
vmem[547] = 8'd105;
vmem[548] = 8'd116;
vmem[549] = 8'd117;
vmem[550] = 8'd114;
vmem[551] = 8'd32;
vmem[552] = 8'd115;
vmem[553] = 8'd105;
vmem[554] = 8'd116;
vmem[555] = 8'd32;
vmem[556] = 8'd97;
vmem[557] = 8'd109;
vmem[558] = 8'd101;
vmem[559] = 8'd116;
vmem[560] = 8'd32;
vmem[561] = 8'd110;
vmem[562] = 8'd105;
vmem[563] = 8'd115;
vmem[564] = 8'd108;
vmem[565] = 8'd32;
vmem[566] = 8'd97;
vmem[567] = 8'd117;
vmem[568] = 8'd103;
vmem[569] = 8'd117;
vmem[570] = 8'd101;
vmem[571] = 8'd46;
vmem[572] = 8'd32;
vmem[573] = 8'd78;
vmem[574] = 8'd117;
vmem[575] = 8'd108;
vmem[576] = 8'd108;
vmem[577] = 8'd97;
vmem[578] = 8'd109;
vmem[579] = 8'd32;
vmem[580] = 8'd118;
vmem[581] = 8'd101;
vmem[582] = 8'd110;
vmem[583] = 8'd101;
vmem[584] = 8'd110;
vmem[585] = 8'd97;
vmem[586] = 8'd116;
vmem[587] = 8'd105;
vmem[588] = 8'd115;
vmem[589] = 8'd32;
vmem[590] = 8'd115;
vmem[591] = 8'd101;
vmem[592] = 8'd109;
vmem[593] = 8'd32;
vmem[594] = 8'd113;
vmem[595] = 8'd117;
vmem[596] = 8'd105;
vmem[597] = 8'd115;
vmem[598] = 8'd32;
vmem[599] = 8'd101;
vmem[600] = 8'd114;
vmem[601] = 8'd97;
vmem[602] = 8'd116;
vmem[603] = 8'd32;
vmem[604] = 8'd102;
vmem[605] = 8'd114;
vmem[606] = 8'd105;
vmem[607] = 8'd110;
vmem[608] = 8'd103;
vmem[609] = 8'd105;
vmem[610] = 8'd108;
vmem[611] = 8'd108;
vmem[612] = 8'd97;
vmem[613] = 8'd32;
vmem[614] = 8'd98;
vmem[615] = 8'd108;
vmem[616] = 8'd97;
vmem[617] = 8'd110;
vmem[618] = 8'd100;
vmem[619] = 8'd105;
vmem[620] = 8'd116;
vmem[621] = 8'd46;
vmem[622] = 8'd32;
vmem[623] = 8'd69;
vmem[624] = 8'd116;
vmem[625] = 8'd105;
vmem[626] = 8'd97;
vmem[627] = 8'd109;
vmem[628] = 8'd32;
vmem[629] = 8'd118;
vmem[630] = 8'd105;
vmem[631] = 8'd118;
vmem[632] = 8'd101;
vmem[633] = 8'd114;
vmem[634] = 8'd114;
vmem[635] = 8'd97;
vmem[636] = 8'd32;
vmem[637] = 8'd108;
vmem[638] = 8'd97;
vmem[639] = 8'd111;
vmem[640] = 8'd114;
vmem[641] = 8'd101;
vmem[642] = 8'd101;
vmem[643] = 8'd116;
vmem[644] = 8'd32;
vmem[645] = 8'd116;
vmem[646] = 8'd111;
vmem[647] = 8'd114;
vmem[648] = 8'd116;
vmem[649] = 8'd111;
vmem[650] = 8'd114;
vmem[651] = 8'd32;
vmem[652] = 8'd110;
vmem[653] = 8'd111;
vmem[654] = 8'd110;
vmem[655] = 8'd32;
vmem[656] = 8'd116;
vmem[657] = 8'd105;
vmem[658] = 8'd110;
vmem[659] = 8'd99;
vmem[660] = 8'd105;
vmem[661] = 8'd100;
vmem[662] = 8'd117;
vmem[663] = 8'd110;
vmem[664] = 8'd116;
vmem[665] = 8'd46;
vmem[666] = 8'd32;
vmem[667] = 8'd86;
vmem[668] = 8'd101;
vmem[669] = 8'd115;
vmem[670] = 8'd116;
vmem[671] = 8'd105;
vmem[672] = 8'd98;
vmem[673] = 8'd117;
vmem[674] = 8'd108;
vmem[675] = 8'd117;
vmem[676] = 8'd109;
vmem[677] = 8'd32;
vmem[678] = 8'd115;
vmem[679] = 8'd105;
vmem[680] = 8'd116;
vmem[681] = 8'd32;
vmem[682] = 8'd97;
vmem[683] = 8'd109;
vmem[684] = 8'd101;
vmem[685] = 8'd116;
vmem[686] = 8'd32;
vmem[687] = 8'd102;
vmem[688] = 8'd105;
vmem[689] = 8'd110;
vmem[690] = 8'd105;
vmem[691] = 8'd98;
vmem[692] = 8'd117;
vmem[693] = 8'd115;
vmem[694] = 8'd32;
vmem[695] = 8'd117;
vmem[696] = 8'd114;
vmem[697] = 8'd110;
vmem[698] = 8'd97;
vmem[699] = 8'd46;
vmem[700] = 8'd32;
vmem[701] = 8'd85;
vmem[702] = 8'd116;
vmem[703] = 8'd32;
vmem[704] = 8'd108;
vmem[705] = 8'd101;
vmem[706] = 8'd99;
vmem[707] = 8'd116;
vmem[708] = 8'd117;
vmem[709] = 8'd115;
vmem[710] = 8'd32;
vmem[711] = 8'd110;
vmem[712] = 8'd117;
vmem[713] = 8'd108;
vmem[714] = 8'd108;
vmem[715] = 8'd97;
vmem[716] = 8'd44;
vmem[717] = 8'd32;
vmem[718] = 8'd99;
vmem[719] = 8'd111;
vmem[720] = 8'd110;
vmem[721] = 8'd118;
vmem[722] = 8'd97;
vmem[723] = 8'd108;
vmem[724] = 8'd108;
vmem[725] = 8'd105;
vmem[726] = 8'd115;
vmem[727] = 8'd32;
vmem[728] = 8'd110;
vmem[729] = 8'd101;
vmem[730] = 8'd99;
vmem[731] = 8'd32;
vmem[732] = 8'd108;
vmem[733] = 8'd117;
vmem[734] = 8'd99;
vmem[735] = 8'd116;
vmem[736] = 8'd117;
vmem[737] = 8'd115;
vmem[738] = 8'd32;
vmem[739] = 8'd110;
vmem[740] = 8'd101;
vmem[741] = 8'd99;
vmem[742] = 8'd44;
vmem[743] = 8'd32;
vmem[744] = 8'd108;
vmem[745] = 8'd97;
vmem[746] = 8'd99;
vmem[747] = 8'd105;
vmem[748] = 8'd110;
vmem[749] = 8'd105;
vmem[750] = 8'd97;
vmem[751] = 8'd32;
vmem[752] = 8'd97;
vmem[753] = 8'd116;
vmem[754] = 8'd32;
vmem[755] = 8'd106;
vmem[756] = 8'd117;
vmem[757] = 8'd115;
vmem[758] = 8'd116;
vmem[759] = 8'd111;
vmem[760] = 8'd46;
vmem[761] = 8'd32;
vmem[762] = 8'd85;
vmem[763] = 8'd116;
vmem[764] = 8'd32;
vmem[765] = 8'd101;
vmem[766] = 8'd114;
vmem[767] = 8'd97;
vmem[768] = 8'd116;
vmem[769] = 8'd32;
vmem[770] = 8'd101;
vmem[771] = 8'd120;
vmem[772] = 8'd44;
vmem[773] = 8'd32;
vmem[774] = 8'd111;
vmem[775] = 8'd114;
vmem[776] = 8'd110;
vmem[777] = 8'd97;
vmem[778] = 8'd114;
vmem[779] = 8'd101;
vmem[780] = 8'd32;
vmem[781] = 8'd101;
vmem[782] = 8'd116;
vmem[783] = 8'd32;
vmem[784] = 8'd101;
vmem[785] = 8'd103;
vmem[786] = 8'd101;
vmem[787] = 8'd115;
vmem[788] = 8'd116;
vmem[789] = 8'd97;
vmem[790] = 8'd115;
vmem[791] = 8'd32;
vmem[792] = 8'd115;
vmem[793] = 8'd105;
vmem[794] = 8'd116;
vmem[795] = 8'd32;
vmem[796] = 8'd97;
vmem[797] = 8'd109;
vmem[798] = 8'd101;
vmem[799] = 8'd116;
vmem[800] = 8'd44;
vmem[801] = 8'd32;
vmem[802] = 8'd115;
vmem[803] = 8'd99;
vmem[804] = 8'd101;
vmem[805] = 8'd108;
vmem[806] = 8'd101;
vmem[807] = 8'd114;
vmem[808] = 8'd105;
vmem[809] = 8'd115;
vmem[810] = 8'd113;
vmem[811] = 8'd117;
vmem[812] = 8'd101;
vmem[813] = 8'd32;
vmem[814] = 8'd101;
vmem[815] = 8'd103;
vmem[816] = 8'd101;
vmem[817] = 8'd116;
vmem[818] = 8'd32;
vmem[819] = 8'd108;
vmem[820] = 8'd105;
vmem[821] = 8'd103;
vmem[822] = 8'd117;
vmem[823] = 8'd108;
vmem[824] = 8'd97;
vmem[825] = 8'd46;
vmem[826] = 8'd32;
vmem[827] = 8'd78;
vmem[828] = 8'd117;
vmem[829] = 8'd108;
vmem[830] = 8'd108;
vmem[831] = 8'd97;
vmem[832] = 8'd32;
vmem[833] = 8'd101;
vmem[834] = 8'd108;
vmem[835] = 8'd101;
vmem[836] = 8'd109;
vmem[837] = 8'd101;
vmem[838] = 8'd110;
vmem[839] = 8'd116;
vmem[840] = 8'd117;
vmem[841] = 8'd109;
vmem[842] = 8'd32;
vmem[843] = 8'd110;
vmem[844] = 8'd105;
vmem[845] = 8'd115;
vmem[846] = 8'd105;
vmem[847] = 8'd32;
vmem[848] = 8'd97;
vmem[849] = 8'd116;
vmem[850] = 8'd32;
vmem[851] = 8'd116;
vmem[852] = 8'd117;
vmem[853] = 8'd114;
vmem[854] = 8'd112;
vmem[855] = 8'd105;
vmem[856] = 8'd115;
vmem[857] = 8'd32;
vmem[858] = 8'd118;
vmem[859] = 8'd101;
vmem[860] = 8'd104;
vmem[861] = 8'd105;
vmem[862] = 8'd99;
vmem[863] = 8'd117;
vmem[864] = 8'd108;
vmem[865] = 8'd97;
vmem[866] = 8'd44;
vmem[867] = 8'd32;
vmem[868] = 8'd110;
vmem[869] = 8'd111;
vmem[870] = 8'd110;
vmem[871] = 8'd32;
vmem[872] = 8'd118;
vmem[873] = 8'd101;
vmem[874] = 8'd104;
vmem[875] = 8'd105;
vmem[876] = 8'd99;
vmem[877] = 8'd117;
vmem[878] = 8'd108;
vmem[879] = 8'd97;
vmem[880] = 8'd32;
vmem[881] = 8'd109;
vmem[882] = 8'd97;
vmem[883] = 8'd115;
vmem[884] = 8'd115;
vmem[885] = 8'd97;
vmem[886] = 8'd32;
vmem[887] = 8'd112;
vmem[888] = 8'd108;
vmem[889] = 8'd97;
vmem[890] = 8'd99;
vmem[891] = 8'd101;
vmem[892] = 8'd114;
vmem[893] = 8'd97;
vmem[894] = 8'd116;
vmem[895] = 8'd46;
vmem[896] = 8'd32;
vmem[897] = 8'd80;
vmem[898] = 8'd104;
vmem[899] = 8'd97;
vmem[900] = 8'd115;
vmem[901] = 8'd101;
vmem[902] = 8'd108;
vmem[903] = 8'd108;
vmem[904] = 8'd117;
vmem[905] = 8'd115;
vmem[906] = 8'd32;
vmem[907] = 8'd99;
vmem[908] = 8'd111;
vmem[909] = 8'd109;
vmem[910] = 8'd109;
vmem[911] = 8'd111;
vmem[912] = 8'd100;
vmem[913] = 8'd111;
vmem[914] = 8'd32;
vmem[915] = 8'd109;
vmem[916] = 8'd101;
vmem[917] = 8'd116;
vmem[918] = 8'd117;
vmem[919] = 8'd115;
vmem[920] = 8'd32;
vmem[921] = 8'd97;
vmem[922] = 8'd116;
vmem[923] = 8'd32;
vmem[924] = 8'd101;
vmem[925] = 8'd114;
vmem[926] = 8'd111;
vmem[927] = 8'd115;
vmem[928] = 8'd32;
vmem[929] = 8'd101;
vmem[930] = 8'd103;
vmem[931] = 8'd101;
vmem[932] = 8'd115;
vmem[933] = 8'd116;
vmem[934] = 8'd97;
vmem[935] = 8'd115;
vmem[936] = 8'd44;
vmem[937] = 8'd32;
vmem[938] = 8'd118;
vmem[939] = 8'd105;
vmem[940] = 8'd116;
vmem[941] = 8'd97;
vmem[942] = 8'd101;
vmem[943] = 8'd32;
vmem[944] = 8'd115;
vmem[945] = 8'd117;
vmem[946] = 8'd115;
vmem[947] = 8'd99;
vmem[948] = 8'd105;
vmem[949] = 8'd112;
vmem[950] = 8'd105;
vmem[951] = 8'd116;
vmem[952] = 8'd32;
vmem[953] = 8'd100;
vmem[954] = 8'd105;
vmem[955] = 8'd97;
vmem[956] = 8'd109;
vmem[957] = 8'd32;
vmem[958] = 8'd105;
vmem[959] = 8'd109;
vmem[960] = 8'd112;
vmem[961] = 8'd101;
vmem[962] = 8'd114;
vmem[963] = 8'd100;
vmem[964] = 8'd105;
vmem[965] = 8'd101;
vmem[966] = 8'd116;
vmem[967] = 8'd46;
vmem[968] = 8'd32;
vmem[969] = 8'd73;
vmem[970] = 8'd110;
vmem[971] = 8'd116;
vmem[972] = 8'd101;
vmem[973] = 8'd103;
vmem[974] = 8'd101;
vmem[975] = 8'd114;
vmem[976] = 8'd32;
vmem[977] = 8'd97;
vmem[978] = 8'd108;
vmem[979] = 8'd105;
vmem[980] = 8'd113;
vmem[981] = 8'd117;
vmem[982] = 8'd101;
vmem[983] = 8'd116;
vmem[984] = 8'd32;
vmem[985] = 8'd97;
vmem[986] = 8'd108;
vmem[987] = 8'd105;
vmem[988] = 8'd113;
vmem[989] = 8'd117;
vmem[990] = 8'd97;
vmem[991] = 8'd109;
vmem[992] = 8'd32;
vmem[993] = 8'd118;
vmem[994] = 8'd101;
vmem[995] = 8'd108;
vmem[996] = 8'd105;
vmem[997] = 8'd116;
vmem[998] = 8'd32;
vmem[999] = 8'd97;
vmem[1000] = 8'd32;
vmem[1001] = 8'd102;
vmem[1002] = 8'd101;
vmem[1003] = 8'd117;
vmem[1004] = 8'd103;
vmem[1005] = 8'd105;
vmem[1006] = 8'd97;
vmem[1007] = 8'd116;
vmem[1008] = 8'd46;
vmem[1009] = 8'd32;
vmem[1010] = 8'd83;
vmem[1011] = 8'd117;
vmem[1012] = 8'd115;
vmem[1013] = 8'd112;
vmem[1014] = 8'd101;
vmem[1015] = 8'd110;
vmem[1016] = 8'd100;
vmem[1017] = 8'd105;
vmem[1018] = 8'd115;
vmem[1019] = 8'd115;
vmem[1020] = 8'd101;
vmem[1021] = 8'd32;
vmem[1022] = 8'd118;
vmem[1023] = 8'd105;
vmem[1024] = 8'd116;
vmem[1025] = 8'd97;
vmem[1026] = 8'd101;
vmem[1027] = 8'd32;
vmem[1028] = 8'd115;
vmem[1029] = 8'd97;
vmem[1030] = 8'd103;
vmem[1031] = 8'd105;
vmem[1032] = 8'd116;
vmem[1033] = 8'd116;
vmem[1034] = 8'd105;
vmem[1035] = 8'd115;
vmem[1036] = 8'd32;
vmem[1037] = 8'd109;
vmem[1038] = 8'd97;
vmem[1039] = 8'd103;
vmem[1040] = 8'd110;
vmem[1041] = 8'd97;
vmem[1042] = 8'd46;
vmem[1043] = 8'd32;
vmem[1044] = 8'd78;
vmem[1045] = 8'd117;
vmem[1046] = 8'd110;
vmem[1047] = 8'd99;
vmem[1048] = 8'd32;
vmem[1049] = 8'd109;
vmem[1050] = 8'd97;
vmem[1051] = 8'd108;
vmem[1052] = 8'd101;
vmem[1053] = 8'd115;
vmem[1054] = 8'd117;
vmem[1055] = 8'd97;
vmem[1056] = 8'd100;
vmem[1057] = 8'd97;
vmem[1058] = 8'd32;
vmem[1059] = 8'd109;
vmem[1060] = 8'd97;
vmem[1061] = 8'd115;
vmem[1062] = 8'd115;
vmem[1063] = 8'd97;
vmem[1064] = 8'd32;
vmem[1065] = 8'd108;
vmem[1066] = 8'd101;
vmem[1067] = 8'd99;
vmem[1068] = 8'd116;
vmem[1069] = 8'd117;
vmem[1070] = 8'd115;
vmem[1071] = 8'd44;
vmem[1072] = 8'd32;
vmem[1073] = 8'd117;
vmem[1074] = 8'd116;
vmem[1075] = 8'd32;
vmem[1076] = 8'd103;
vmem[1077] = 8'd114;
vmem[1078] = 8'd97;
vmem[1079] = 8'd118;
vmem[1080] = 8'd105;
vmem[1081] = 8'd100;
vmem[1082] = 8'd97;
vmem[1083] = 8'd32;
vmem[1084] = 8'd100;
vmem[1085] = 8'd111;
vmem[1086] = 8'd108;
vmem[1087] = 8'd111;
vmem[1088] = 8'd114;
vmem[1089] = 8'd32;
vmem[1090] = 8'd105;
vmem[1091] = 8'd110;
vmem[1092] = 8'd116;
vmem[1093] = 8'd101;
vmem[1094] = 8'd114;
vmem[1095] = 8'd100;
vmem[1096] = 8'd117;
vmem[1097] = 8'd109;
vmem[1098] = 8'd32;
vmem[1099] = 8'd115;
vmem[1100] = 8'd101;
vmem[1101] = 8'd100;
vmem[1102] = 8'd46;
vmem[1103] = 8'd32;
vmem[1104] = 8'd70;
vmem[1105] = 8'd117;
vmem[1106] = 8'd115;
vmem[1107] = 8'd99;
vmem[1108] = 8'd101;
vmem[1109] = 8'd32;
vmem[1110] = 8'd109;
vmem[1111] = 8'd97;
vmem[1112] = 8'd116;
vmem[1113] = 8'd116;
vmem[1114] = 8'd105;
vmem[1115] = 8'd115;
vmem[1116] = 8'd32;
vmem[1117] = 8'd109;
vmem[1118] = 8'd105;
vmem[1119] = 8'd32;
vmem[1120] = 8'd118;
vmem[1121] = 8'd101;
vmem[1122] = 8'd108;
vmem[1123] = 8'd32;
vmem[1124] = 8'd115;
vmem[1125] = 8'd97;
vmem[1126] = 8'd112;
vmem[1127] = 8'd105;
vmem[1128] = 8'd101;
vmem[1129] = 8'd110;
vmem[1130] = 8'd32;
vmem[1131] = 8'd105;
vmem[1132] = 8'd109;
vmem[1133] = 8'd112;
vmem[1134] = 8'd101;
vmem[1135] = 8'd114;
vmem[1136] = 8'd100;
vmem[1137] = 8'd105;
vmem[1138] = 8'd101;
vmem[1139] = 8'd116;
vmem[1140] = 8'd44;
vmem[1141] = 8'd32;
vmem[1142] = 8'd101;
vmem[1143] = 8'd117;
vmem[1144] = 8'd105;
vmem[1145] = 8'd115;
vmem[1146] = 8'd109;
vmem[1147] = 8'd111;
vmem[1148] = 8'd100;
vmem[1149] = 8'd32;
vmem[1150] = 8'd102;
vmem[1151] = 8'd114;
vmem[1152] = 8'd105;
vmem[1153] = 8'd110;
vmem[1154] = 8'd103;
vmem[1155] = 8'd105;
vmem[1156] = 8'd108;
vmem[1157] = 8'd108;
vmem[1158] = 8'd97;
vmem[1159] = 8'd32;
vmem[1160] = 8'd101;
vmem[1161] = 8'd110;
vmem[1162] = 8'd105;
vmem[1163] = 8'd109;
vmem[1164] = 8'd32;
vmem[1165] = 8'd108;
vmem[1166] = 8'd97;
vmem[1167] = 8'd111;
vmem[1168] = 8'd114;
vmem[1169] = 8'd101;
vmem[1170] = 8'd101;
vmem[1171] = 8'd116;
vmem[1172] = 8'd46;
vmem[1173] = 8'd32;
vmem[1174] = 8'd68;
vmem[1175] = 8'd111;
vmem[1176] = 8'd110;
vmem[1177] = 8'd101;
vmem[1178] = 8'd99;
vmem[1179] = 8'd32;
vmem[1180] = 8'd118;
vmem[1181] = 8'd111;
vmem[1182] = 8'd108;
vmem[1183] = 8'd117;
vmem[1184] = 8'd116;
vmem[1185] = 8'd112;
vmem[1186] = 8'd97;
vmem[1187] = 8'd116;
vmem[1188] = 8'd44;
vmem[1189] = 8'd32;
vmem[1190] = 8'd116;
vmem[1191] = 8'd117;
vmem[1192] = 8'd114;
vmem[1193] = 8'd112;
vmem[1194] = 8'd105;
vmem[1195] = 8'd115;
vmem[1196] = 8'd32;
vmem[1197] = 8'd97;
vmem[1198] = 8'd99;
vmem[1199] = 8'd32;
vmem[1200] = 8'd118;
vmem[1201] = 8'd101;
vmem[1202] = 8'd104;
vmem[1203] = 8'd105;
vmem[1204] = 8'd99;
vmem[1205] = 8'd117;
vmem[1206] = 8'd108;
vmem[1207] = 8'd97;
vmem[1208] = 8'd32;
vmem[1209] = 8'd104;
vmem[1210] = 8'd101;
vmem[1211] = 8'd110;
vmem[1212] = 8'd100;
vmem[1213] = 8'd114;
vmem[1214] = 8'd101;
vmem[1215] = 8'd114;
vmem[1216] = 8'd105;
vmem[1217] = 8'd116;
vmem[1218] = 8'd44;
vmem[1219] = 8'd32;
vmem[1220] = 8'd111;
vmem[1221] = 8'd100;
vmem[1222] = 8'd105;
vmem[1223] = 8'd111;
vmem[1224] = 8'd32;
vmem[1225] = 8'd115;
vmem[1226] = 8'd97;
vmem[1227] = 8'd112;
vmem[1228] = 8'd105;
vmem[1229] = 8'd101;
vmem[1230] = 8'd110;
vmem[1231] = 8'd32;
vmem[1232] = 8'd112;
vmem[1233] = 8'd104;
vmem[1234] = 8'd97;
vmem[1235] = 8'd114;
vmem[1236] = 8'd101;
vmem[1237] = 8'd116;
vmem[1238] = 8'd114;
vmem[1239] = 8'd97;
vmem[1240] = 8'd32;
vmem[1241] = 8'd115;
vmem[1242] = 8'd101;
vmem[1243] = 8'd109;
vmem[1244] = 8'd44;
vmem[1245] = 8'd32;
vmem[1246] = 8'd117;
vmem[1247] = 8'd116;
vmem[1248] = 8'd32;
vmem[1249] = 8'd109;
vmem[1250] = 8'd97;
vmem[1251] = 8'd120;
vmem[1252] = 8'd105;
vmem[1253] = 8'd109;
vmem[1254] = 8'd117;
vmem[1255] = 8'd115;
vmem[1256] = 8'd32;
vmem[1257] = 8'd109;
vmem[1258] = 8'd97;
vmem[1259] = 8'd103;
vmem[1260] = 8'd110;
vmem[1261] = 8'd97;
vmem[1262] = 8'd32;
vmem[1263] = 8'd112;
vmem[1264] = 8'd117;
vmem[1265] = 8'd114;
vmem[1266] = 8'd117;
vmem[1267] = 8'd115;
vmem[1268] = 8'd32;
vmem[1269] = 8'd97;
vmem[1270] = 8'd99;
vmem[1271] = 8'd32;
vmem[1272] = 8'd111;
vmem[1273] = 8'd100;
vmem[1274] = 8'd105;
vmem[1275] = 8'd111;
vmem[1276] = 8'd46;
vmem[1277] = 8'd32;
vmem[1278] = 8'd78;
vmem[1279] = 8'd117;
vmem[1280] = 8'd108;
vmem[1281] = 8'd108;
vmem[1282] = 8'd97;
vmem[1283] = 8'd32;
vmem[1284] = 8'd118;
vmem[1285] = 8'd105;
vmem[1286] = 8'd116;
vmem[1287] = 8'd97;
vmem[1288] = 8'd101;
vmem[1289] = 8'd32;
vmem[1290] = 8'd116;
vmem[1291] = 8'd117;
vmem[1292] = 8'd114;
vmem[1293] = 8'd112;
vmem[1294] = 8'd105;
vmem[1295] = 8'd115;
vmem[1296] = 8'd32;
vmem[1297] = 8'd100;
vmem[1298] = 8'd105;
vmem[1299] = 8'd103;
vmem[1300] = 8'd110;
vmem[1301] = 8'd105;
vmem[1302] = 8'd115;
vmem[1303] = 8'd115;
vmem[1304] = 8'd105;
vmem[1305] = 8'd109;
vmem[1306] = 8'd44;
vmem[1307] = 8'd32;
vmem[1308] = 8'd97;
vmem[1309] = 8'd108;
vmem[1310] = 8'd105;
vmem[1311] = 8'd113;
vmem[1312] = 8'd117;
vmem[1313] = 8'd97;
vmem[1314] = 8'd109;
vmem[1315] = 8'd32;
vmem[1316] = 8'd101;
vmem[1317] = 8'd114;
vmem[1318] = 8'd111;
vmem[1319] = 8'd115;
vmem[1320] = 8'd32;
vmem[1321] = 8'd101;
vmem[1322] = 8'd117;
vmem[1323] = 8'd44;
vmem[1324] = 8'd32;
vmem[1325] = 8'd102;
vmem[1326] = 8'd114;
vmem[1327] = 8'd105;
vmem[1328] = 8'd110;
vmem[1329] = 8'd103;
vmem[1330] = 8'd105;
vmem[1331] = 8'd108;
vmem[1332] = 8'd108;
vmem[1333] = 8'd97;
vmem[1334] = 8'd32;
vmem[1335] = 8'd109;
vmem[1336] = 8'd97;
vmem[1337] = 8'd115;
vmem[1338] = 8'd115;
vmem[1339] = 8'd97;
vmem[1340] = 8'd46;
vmem[1341] = 8'd32;
vmem[1342] = 8'd78;
vmem[1343] = 8'd97;
vmem[1344] = 8'd109;
vmem[1345] = 8'd32;
vmem[1346] = 8'd99;
vmem[1347] = 8'd111;
vmem[1348] = 8'd110;
vmem[1349] = 8'd115;
vmem[1350] = 8'd101;
vmem[1351] = 8'd99;
vmem[1352] = 8'd116;
vmem[1353] = 8'd101;
vmem[1354] = 8'd116;
vmem[1355] = 8'd117;
vmem[1356] = 8'd114;
vmem[1357] = 8'd32;
vmem[1358] = 8'd110;
vmem[1359] = 8'd105;
vmem[1360] = 8'd115;
vmem[1361] = 8'd108;
vmem[1362] = 8'd32;
vmem[1363] = 8'd105;
vmem[1364] = 8'd100;
vmem[1365] = 8'd32;
vmem[1366] = 8'd100;
vmem[1367] = 8'd111;
vmem[1368] = 8'd108;
vmem[1369] = 8'd111;
vmem[1370] = 8'd114;
vmem[1371] = 8'd32;
vmem[1372] = 8'd99;
vmem[1373] = 8'd111;
vmem[1374] = 8'd110;
vmem[1375] = 8'd118;
vmem[1376] = 8'd97;
vmem[1377] = 8'd108;
vmem[1378] = 8'd108;
vmem[1379] = 8'd105;
vmem[1380] = 8'd115;
vmem[1381] = 8'd32;
vmem[1382] = 8'd100;
vmem[1383] = 8'd105;
vmem[1384] = 8'd103;
vmem[1385] = 8'd110;
vmem[1386] = 8'd105;
vmem[1387] = 8'd115;
vmem[1388] = 8'd115;
vmem[1389] = 8'd105;
vmem[1390] = 8'd109;
vmem[1391] = 8'd46;
vmem[1392] = 8'd32;
vmem[1393] = 8'd81;
vmem[1394] = 8'd117;
vmem[1395] = 8'd105;
vmem[1396] = 8'd115;
vmem[1397] = 8'd113;
vmem[1398] = 8'd117;
vmem[1399] = 8'd101;
vmem[1400] = 8'd32;
vmem[1401] = 8'd115;
vmem[1402] = 8'd117;
vmem[1403] = 8'd115;
vmem[1404] = 8'd99;
vmem[1405] = 8'd105;
vmem[1406] = 8'd112;
vmem[1407] = 8'd105;
vmem[1408] = 8'd116;
vmem[1409] = 8'd32;
vmem[1410] = 8'd112;
vmem[1411] = 8'd111;
vmem[1412] = 8'd114;
vmem[1413] = 8'd116;
vmem[1414] = 8'd116;
vmem[1415] = 8'd105;
vmem[1416] = 8'd116;
vmem[1417] = 8'd111;
vmem[1418] = 8'd114;
vmem[1419] = 8'd32;
vmem[1420] = 8'd100;
vmem[1421] = 8'd117;
vmem[1422] = 8'd105;
vmem[1423] = 8'd32;
vmem[1424] = 8'd105;
vmem[1425] = 8'd100;
vmem[1426] = 8'd32;
vmem[1427] = 8'd99;
vmem[1428] = 8'd111;
vmem[1429] = 8'd110;
vmem[1430] = 8'd103;
vmem[1431] = 8'd117;
vmem[1432] = 8'd101;
vmem[1433] = 8'd46;
vmem[1434] = 8'd32;
vmem[1435] = 8'd85;
vmem[1436] = 8'd116;
vmem[1437] = 8'd32;
vmem[1438] = 8'd102;
vmem[1439] = 8'd114;
vmem[1440] = 8'd105;
vmem[1441] = 8'd110;
vmem[1442] = 8'd103;
vmem[1443] = 8'd105;
vmem[1444] = 8'd108;
vmem[1445] = 8'd108;
vmem[1446] = 8'd97;
vmem[1447] = 8'd32;
vmem[1448] = 8'd101;
vmem[1449] = 8'd103;
vmem[1450] = 8'd101;
vmem[1451] = 8'd116;
vmem[1452] = 8'd32;
vmem[1453] = 8'd114;
vmem[1454] = 8'd105;
vmem[1455] = 8'd115;
vmem[1456] = 8'd117;
vmem[1457] = 8'd115;
vmem[1458] = 8'd32;
vmem[1459] = 8'd118;
vmem[1460] = 8'd101;
vmem[1461] = 8'd108;
vmem[1462] = 8'd32;
vmem[1463] = 8'd115;
vmem[1464] = 8'd97;
vmem[1465] = 8'd103;
vmem[1466] = 8'd105;
vmem[1467] = 8'd116;
vmem[1468] = 8'd116;
vmem[1469] = 8'd105;
vmem[1470] = 8'd115;
vmem[1471] = 8'd46;
vmem[1472] = 8'd32;
vmem[1473] = 8'd77;
vmem[1474] = 8'd97;
vmem[1475] = 8'd101;
vmem[1476] = 8'd99;
vmem[1477] = 8'd101;
vmem[1478] = 8'd110;
vmem[1479] = 8'd97;
vmem[1480] = 8'd115;
vmem[1481] = 8'd32;
vmem[1482] = 8'd105;
vmem[1483] = 8'd110;
vmem[1484] = 8'd116;
vmem[1485] = 8'd101;
vmem[1486] = 8'd114;
vmem[1487] = 8'd100;
vmem[1488] = 8'd117;
vmem[1489] = 8'd109;
vmem[1490] = 8'd32;
vmem[1491] = 8'd118;
vmem[1492] = 8'd101;
vmem[1493] = 8'd108;
vmem[1494] = 8'd105;
vmem[1495] = 8'd116;
vmem[1496] = 8'd32;
vmem[1497] = 8'd110;
vmem[1498] = 8'd111;
vmem[1499] = 8'd110;
vmem[1500] = 8'd32;
vmem[1501] = 8'd102;
vmem[1502] = 8'd97;
vmem[1503] = 8'd117;
vmem[1504] = 8'd99;
vmem[1505] = 8'd105;
vmem[1506] = 8'd98;
vmem[1507] = 8'd117;
vmem[1508] = 8'd115;
vmem[1509] = 8'd32;
vmem[1510] = 8'd109;
vmem[1511] = 8'd97;
vmem[1512] = 8'd120;
vmem[1513] = 8'd105;
vmem[1514] = 8'd109;
vmem[1515] = 8'd117;
vmem[1516] = 8'd115;
vmem[1517] = 8'd46;
vmem[1518] = 8'd32;
vmem[1519] = 8'd78;
vmem[1520] = 8'd117;
vmem[1521] = 8'd110;
vmem[1522] = 8'd99;
vmem[1523] = 8'd32;
vmem[1524] = 8'd110;
vmem[1525] = 8'd101;
vmem[1526] = 8'd99;
vmem[1527] = 8'd32;
vmem[1528] = 8'd115;
vmem[1529] = 8'd97;
vmem[1530] = 8'd103;
vmem[1531] = 8'd105;
vmem[1532] = 8'd116;
vmem[1533] = 8'd116;
vmem[1534] = 8'd105;
vmem[1535] = 8'd115;
vmem[1536] = 8'd32;
vmem[1537] = 8'd114;
vmem[1538] = 8'd105;
vmem[1539] = 8'd115;
vmem[1540] = 8'd117;
vmem[1541] = 8'd115;
vmem[1542] = 8'd44;
vmem[1543] = 8'd32;
vmem[1544] = 8'd97;
vmem[1545] = 8'd108;
vmem[1546] = 8'd105;
vmem[1547] = 8'd113;
vmem[1548] = 8'd117;
vmem[1549] = 8'd97;
vmem[1550] = 8'd109;
vmem[1551] = 8'd32;
vmem[1552] = 8'd116;
vmem[1553] = 8'd101;
vmem[1554] = 8'd109;
vmem[1555] = 8'd112;
vmem[1556] = 8'd111;
vmem[1557] = 8'd114;
vmem[1558] = 8'd32;
vmem[1559] = 8'd109;
vmem[1560] = 8'd105;
vmem[1561] = 8'd46;
vmem[1562] = 8'd32;
vmem[1563] = 8'd78;
vmem[1564] = 8'd117;
vmem[1565] = 8'd108;
vmem[1566] = 8'd108;
vmem[1567] = 8'd97;
vmem[1568] = 8'd109;
vmem[1569] = 8'd32;
vmem[1570] = 8'd110;
vmem[1571] = 8'd105;
vmem[1572] = 8'd115;
vmem[1573] = 8'd105;
vmem[1574] = 8'd32;
vmem[1575] = 8'd97;
vmem[1576] = 8'd114;
vmem[1577] = 8'd99;
vmem[1578] = 8'd117;
vmem[1579] = 8'd44;
vmem[1580] = 8'd32;
vmem[1581] = 8'd102;
vmem[1582] = 8'd97;
vmem[1583] = 8'd117;
vmem[1584] = 8'd99;
vmem[1585] = 8'd105;
vmem[1586] = 8'd98;
vmem[1587] = 8'd117;
vmem[1588] = 8'd115;
vmem[1589] = 8'd32;
vmem[1590] = 8'd117;
vmem[1591] = 8'd116;
vmem[1592] = 8'd32;
vmem[1593] = 8'd109;
vmem[1594] = 8'd97;
vmem[1595] = 8'd117;
vmem[1596] = 8'd114;
vmem[1597] = 8'd105;
vmem[1598] = 8'd115;
vmem[1599] = 8'd32;
vmem[1600] = 8'd116;
vmem[1601] = 8'd101;
vmem[1602] = 8'd109;
vmem[1603] = 8'd112;
vmem[1604] = 8'd117;
vmem[1605] = 8'd115;
vmem[1606] = 8'd44;
vmem[1607] = 8'd32;
vmem[1608] = 8'd118;
vmem[1609] = 8'd101;
vmem[1610] = 8'd104;
vmem[1611] = 8'd105;
vmem[1612] = 8'd99;
vmem[1613] = 8'd117;
vmem[1614] = 8'd108;
vmem[1615] = 8'd97;
vmem[1616] = 8'd32;
vmem[1617] = 8'd118;
vmem[1618] = 8'd117;
vmem[1619] = 8'd108;
vmem[1620] = 8'd112;
vmem[1621] = 8'd117;
vmem[1622] = 8'd116;
vmem[1623] = 8'd97;
vmem[1624] = 8'd116;
vmem[1625] = 8'd101;
vmem[1626] = 8'd32;
vmem[1627] = 8'd109;
vmem[1628] = 8'd97;
vmem[1629] = 8'd115;
vmem[1630] = 8'd115;
vmem[1631] = 8'd97;
vmem[1632] = 8'd46;
vmem[1633] = 8'd32;
vmem[1634] = 8'd77;
vmem[1635] = 8'd97;
vmem[1636] = 8'd117;
vmem[1637] = 8'd114;
vmem[1638] = 8'd105;
vmem[1639] = 8'd115;
vmem[1640] = 8'd32;
vmem[1641] = 8'd118;
vmem[1642] = 8'd111;
vmem[1643] = 8'd108;
vmem[1644] = 8'd117;
vmem[1645] = 8'd116;
vmem[1646] = 8'd112;
vmem[1647] = 8'd97;
vmem[1648] = 8'd116;
vmem[1649] = 8'd44;
vmem[1650] = 8'd32;
vmem[1651] = 8'd110;
vmem[1652] = 8'd105;
vmem[1653] = 8'd115;
vmem[1654] = 8'd108;
vmem[1655] = 8'd32;
vmem[1656] = 8'd105;
vmem[1657] = 8'd100;
vmem[1658] = 8'd32;
vmem[1659] = 8'd118;
vmem[1660] = 8'd111;
vmem[1661] = 8'd108;
vmem[1662] = 8'd117;
vmem[1663] = 8'd116;
vmem[1664] = 8'd112;
vmem[1665] = 8'd97;
vmem[1666] = 8'd116;
vmem[1667] = 8'd32;
vmem[1668] = 8'd99;
vmem[1669] = 8'd111;
vmem[1670] = 8'd109;
vmem[1671] = 8'd109;
vmem[1672] = 8'd111;
vmem[1673] = 8'd100;
vmem[1674] = 8'd111;
vmem[1675] = 8'd44;
vmem[1676] = 8'd32;
vmem[1677] = 8'd101;
vmem[1678] = 8'd120;
vmem[1679] = 8'd32;
vmem[1680] = 8'd115;
vmem[1681] = 8'd101;
vmem[1682] = 8'd109;
vmem[1683] = 8'd32;
vmem[1684] = 8'd102;
vmem[1685] = 8'd101;
vmem[1686] = 8'd117;
vmem[1687] = 8'd103;
vmem[1688] = 8'd105;
vmem[1689] = 8'd97;
vmem[1690] = 8'd116;
vmem[1691] = 8'd32;
vmem[1692] = 8'd113;
vmem[1693] = 8'd117;
vmem[1694] = 8'd97;
vmem[1695] = 8'd109;
vmem[1696] = 8'd44;
vmem[1697] = 8'd32;
vmem[1698] = 8'd101;
vmem[1699] = 8'd103;
vmem[1700] = 8'd101;
vmem[1701] = 8'd116;
vmem[1702] = 8'd32;
vmem[1703] = 8'd112;
vmem[1704] = 8'd114;
vmem[1705] = 8'd101;
vmem[1706] = 8'd116;
vmem[1707] = 8'd105;
vmem[1708] = 8'd117;
vmem[1709] = 8'd109;
vmem[1710] = 8'd32;
vmem[1711] = 8'd112;
vmem[1712] = 8'd117;
vmem[1713] = 8'd114;
vmem[1714] = 8'd117;
vmem[1715] = 8'd115;
vmem[1716] = 8'd32;
vmem[1717] = 8'd108;
vmem[1718] = 8'd101;
vmem[1719] = 8'd111;
vmem[1720] = 8'd32;
vmem[1721] = 8'd109;
vmem[1722] = 8'd97;
vmem[1723] = 8'd108;
vmem[1724] = 8'd101;
vmem[1725] = 8'd115;
vmem[1726] = 8'd117;
vmem[1727] = 8'd97;
vmem[1728] = 8'd100;
vmem[1729] = 8'd97;
vmem[1730] = 8'd32;
vmem[1731] = 8'd100;
vmem[1732] = 8'd111;
vmem[1733] = 8'd108;
vmem[1734] = 8'd111;
vmem[1735] = 8'd114;
vmem[1736] = 8'd46;
vmem[1737] = 8'd32;
vmem[1738] = 8'd80;
vmem[1739] = 8'd104;
vmem[1740] = 8'd97;
vmem[1741] = 8'd115;
vmem[1742] = 8'd101;
vmem[1743] = 8'd108;
vmem[1744] = 8'd108;
vmem[1745] = 8'd117;
vmem[1746] = 8'd115;
vmem[1747] = 8'd32;
vmem[1748] = 8'd110;
vmem[1749] = 8'd111;
vmem[1750] = 8'd110;
vmem[1751] = 8'd32;
vmem[1752] = 8'd110;
vmem[1753] = 8'd117;
vmem[1754] = 8'd108;
vmem[1755] = 8'd108;
vmem[1756] = 8'd97;
vmem[1757] = 8'd32;
vmem[1758] = 8'd112;
vmem[1759] = 8'd101;
vmem[1760] = 8'd108;
vmem[1761] = 8'd108;
vmem[1762] = 8'd101;
vmem[1763] = 8'd110;
vmem[1764] = 8'd116;
vmem[1765] = 8'd101;
vmem[1766] = 8'd115;
vmem[1767] = 8'd113;
vmem[1768] = 8'd117;
vmem[1769] = 8'd101;
vmem[1770] = 8'd44;
vmem[1771] = 8'd32;
vmem[1772] = 8'd115;
vmem[1773] = 8'd111;
vmem[1774] = 8'd108;
vmem[1775] = 8'd108;
vmem[1776] = 8'd105;
vmem[1777] = 8'd99;
vmem[1778] = 8'd105;
vmem[1779] = 8'd116;
vmem[1780] = 8'd117;
vmem[1781] = 8'd100;
vmem[1782] = 8'd105;
vmem[1783] = 8'd110;
vmem[1784] = 8'd32;
vmem[1785] = 8'd115;
vmem[1786] = 8'd97;
vmem[1787] = 8'd112;
vmem[1788] = 8'd105;
vmem[1789] = 8'd101;
vmem[1790] = 8'd110;
vmem[1791] = 8'd32;
vmem[1792] = 8'd118;
vmem[1793] = 8'd105;
vmem[1794] = 8'd116;
vmem[1795] = 8'd97;
vmem[1796] = 8'd101;
vmem[1797] = 8'd44;
vmem[1798] = 8'd32;
vmem[1799] = 8'd115;
vmem[1800] = 8'd97;
vmem[1801] = 8'd103;
vmem[1802] = 8'd105;
vmem[1803] = 8'd116;
vmem[1804] = 8'd116;
vmem[1805] = 8'd105;
vmem[1806] = 8'd115;
vmem[1807] = 8'd32;
vmem[1808] = 8'd108;
vmem[1809] = 8'd111;
vmem[1810] = 8'd114;
vmem[1811] = 8'd101;
vmem[1812] = 8'd109;
vmem[1813] = 8'd46;
vmem[1814] = 8'd32;
vmem[1815] = 8'd69;
vmem[1816] = 8'd116;
vmem[1817] = 8'd105;
vmem[1818] = 8'd97;
vmem[1819] = 8'd109;
vmem[1820] = 8'd32;
vmem[1821] = 8'd110;
vmem[1822] = 8'd101;
vmem[1823] = 8'd99;
vmem[1824] = 8'd32;
vmem[1825] = 8'd99;
vmem[1826] = 8'd111;
vmem[1827] = 8'd110;
vmem[1828] = 8'd118;
vmem[1829] = 8'd97;
vmem[1830] = 8'd108;
vmem[1831] = 8'd108;
vmem[1832] = 8'd105;
vmem[1833] = 8'd115;
vmem[1834] = 8'd32;
vmem[1835] = 8'd109;
vmem[1836] = 8'd105;
vmem[1837] = 8'd44;
vmem[1838] = 8'd32;
vmem[1839] = 8'd97;
vmem[1840] = 8'd116;
vmem[1841] = 8'd32;
vmem[1842] = 8'd118;
vmem[1843] = 8'd97;
vmem[1844] = 8'd114;
vmem[1845] = 8'd105;
vmem[1846] = 8'd117;
vmem[1847] = 8'd115;
vmem[1848] = 8'd32;
vmem[1849] = 8'd108;
vmem[1850] = 8'd111;
vmem[1851] = 8'd114;
vmem[1852] = 8'd101;
vmem[1853] = 8'd109;
vmem[1854] = 8'd46;
vmem[1855] = 8'd32;
vmem[1856] = 8'd80;
vmem[1857] = 8'd114;
vmem[1858] = 8'd111;
vmem[1859] = 8'd105;
vmem[1860] = 8'd110;
vmem[1861] = 8'd32;
vmem[1862] = 8'd109;
vmem[1863] = 8'd111;
vmem[1864] = 8'd108;
vmem[1865] = 8'd101;
vmem[1866] = 8'd115;
vmem[1867] = 8'd116;
vmem[1868] = 8'd105;
vmem[1869] = 8'd101;
vmem[1870] = 8'd32;
vmem[1871] = 8'd101;
vmem[1872] = 8'd110;
vmem[1873] = 8'd105;
vmem[1874] = 8'd109;
vmem[1875] = 8'd32;
vmem[1876] = 8'd116;
vmem[1877] = 8'd111;
vmem[1878] = 8'd114;
vmem[1879] = 8'd116;
vmem[1880] = 8'd111;
vmem[1881] = 8'd114;
vmem[1882] = 8'd44;
vmem[1883] = 8'd32;
vmem[1884] = 8'd115;
vmem[1885] = 8'd101;
vmem[1886] = 8'd100;
vmem[1887] = 8'd32;
vmem[1888] = 8'd108;
vmem[1889] = 8'd117;
vmem[1890] = 8'd99;
vmem[1891] = 8'd116;
vmem[1892] = 8'd117;
vmem[1893] = 8'd115;
vmem[1894] = 8'd32;
vmem[1895] = 8'd116;
vmem[1896] = 8'd101;
vmem[1897] = 8'd108;
vmem[1898] = 8'd108;
vmem[1899] = 8'd117;
vmem[1900] = 8'd115;
vmem[1901] = 8'd32;
vmem[1902] = 8'd97;
vmem[1903] = 8'd108;
vmem[1904] = 8'd105;
vmem[1905] = 8'd113;
vmem[1906] = 8'd117;
vmem[1907] = 8'd97;
vmem[1908] = 8'd109;
vmem[1909] = 8'd32;
vmem[1910] = 8'd118;
vmem[1911] = 8'd105;
vmem[1912] = 8'd116;
vmem[1913] = 8'd97;
vmem[1914] = 8'd101;
vmem[1915] = 8'd46;
vmem[1916] = 8'd32;
vmem[1917] = 8'd83;
vmem[1918] = 8'd101;
vmem[1919] = 8'd100;
vmem[1920] = 8'd32;
vmem[1921] = 8'd97;
vmem[1922] = 8'd108;
vmem[1923] = 8'd105;
vmem[1924] = 8'd113;
vmem[1925] = 8'd117;
vmem[1926] = 8'd97;
vmem[1927] = 8'd109;
vmem[1928] = 8'd32;
vmem[1929] = 8'd118;
vmem[1930] = 8'd101;
vmem[1931] = 8'd108;
vmem[1932] = 8'd32;
vmem[1933] = 8'd101;
vmem[1934] = 8'd108;
vmem[1935] = 8'd105;
vmem[1936] = 8'd116;
vmem[1937] = 8'd32;
vmem[1938] = 8'd116;
vmem[1939] = 8'd105;
vmem[1940] = 8'd110;
vmem[1941] = 8'd99;
vmem[1942] = 8'd105;
vmem[1943] = 8'd100;
vmem[1944] = 8'd117;
vmem[1945] = 8'd110;
vmem[1946] = 8'd116;
vmem[1947] = 8'd32;
vmem[1948] = 8'd102;
vmem[1949] = 8'd114;
vmem[1950] = 8'd105;
vmem[1951] = 8'd110;
vmem[1952] = 8'd103;
vmem[1953] = 8'd105;
vmem[1954] = 8'd108;
vmem[1955] = 8'd108;
vmem[1956] = 8'd97;
vmem[1957] = 8'd46;
vmem[1958] = 8'd32;
vmem[1959] = 8'd65;
vmem[1960] = 8'd101;
vmem[1961] = 8'd110;
vmem[1962] = 8'd101;
vmem[1963] = 8'd97;
vmem[1964] = 8'd110;
vmem[1965] = 8'd32;
vmem[1966] = 8'd110;
vmem[1967] = 8'd105;
vmem[1968] = 8'd115;
vmem[1969] = 8'd108;
vmem[1970] = 8'd32;
vmem[1971] = 8'd108;
vmem[1972] = 8'd105;
vmem[1973] = 8'd103;
vmem[1974] = 8'd117;
vmem[1975] = 8'd108;
vmem[1976] = 8'd97;
vmem[1977] = 8'd44;
vmem[1978] = 8'd32;
vmem[1979] = 8'd115;
vmem[1980] = 8'd117;
vmem[1981] = 8'd115;
vmem[1982] = 8'd99;
vmem[1983] = 8'd105;
vmem[1984] = 8'd112;
vmem[1985] = 8'd105;
vmem[1986] = 8'd116;
vmem[1987] = 8'd32;
vmem[1988] = 8'd97;
vmem[1989] = 8'd116;
vmem[1990] = 8'd32;
vmem[1991] = 8'd101;
vmem[1992] = 8'd103;
vmem[1993] = 8'd101;
vmem[1994] = 8'd115;
vmem[1995] = 8'd116;
vmem[1996] = 8'd97;
vmem[1997] = 8'd115;
vmem[1998] = 8'd32;
vmem[1999] = 8'd110;
vmem[2000] = 8'd101;
vmem[2001] = 8'd99;
vmem[2002] = 8'd44;
vmem[2003] = 8'd32;
vmem[2004] = 8'd99;
vmem[2005] = 8'd111;
vmem[2006] = 8'd109;
vmem[2007] = 8'd109;
vmem[2008] = 8'd111;
vmem[2009] = 8'd100;
vmem[2010] = 8'd111;
vmem[2011] = 8'd32;
vmem[2012] = 8'd101;
vmem[2013] = 8'd117;
vmem[2014] = 8'd32;
vmem[2015] = 8'd111;
vmem[2016] = 8'd100;
vmem[2017] = 8'd105;
vmem[2018] = 8'd111;
vmem[2019] = 8'd46;
vmem[2020] = 8'd32;
vmem[2021] = 8'd80;
vmem[2022] = 8'd114;
vmem[2023] = 8'd97;
vmem[2024] = 8'd101;
vmem[2025] = 8'd115;
vmem[2026] = 8'd101;
vmem[2027] = 8'd110;
vmem[2028] = 8'd116;
vmem[2029] = 8'd32;
vmem[2030] = 8'd116;
vmem[2031] = 8'd114;
vmem[2032] = 8'd105;
vmem[2033] = 8'd115;
vmem[2034] = 8'd116;
vmem[2035] = 8'd105;
vmem[2036] = 8'd113;
vmem[2037] = 8'd117;
vmem[2038] = 8'd101;
vmem[2039] = 8'd32;
vmem[2040] = 8'd105;
vmem[2041] = 8'd100;
vmem[2042] = 8'd32;
vmem[2043] = 8'd100;
vmem[2044] = 8'd105;
vmem[2045] = 8'd97;
vmem[2046] = 8'd109;
vmem[2047] = 8'd32;
vmem[2048] = 8'd97;
vmem[2049] = 8'd32;
vmem[2050] = 8'd97;
vmem[2051] = 8'd99;
vmem[2052] = 8'd99;
vmem[2053] = 8'd117;
vmem[2054] = 8'd109;
vmem[2055] = 8'd115;
vmem[2056] = 8'd97;
vmem[2057] = 8'd110;
vmem[2058] = 8'd46;
vmem[2059] = 8'd32;
vmem[2060] = 8'd83;
vmem[2061] = 8'd117;
vmem[2062] = 8'd115;
vmem[2063] = 8'd112;
vmem[2064] = 8'd101;
vmem[2065] = 8'd110;
vmem[2066] = 8'd100;
vmem[2067] = 8'd105;
vmem[2068] = 8'd115;
vmem[2069] = 8'd115;
vmem[2070] = 8'd101;
vmem[2071] = 8'd32;
vmem[2072] = 8'd98;
vmem[2073] = 8'd105;
vmem[2074] = 8'd98;
vmem[2075] = 8'd101;
vmem[2076] = 8'd110;
vmem[2077] = 8'd100;
vmem[2078] = 8'd117;
vmem[2079] = 8'd109;
vmem[2080] = 8'd32;
vmem[2081] = 8'd108;
vmem[2082] = 8'd111;
vmem[2083] = 8'd98;
vmem[2084] = 8'd111;
vmem[2085] = 8'd114;
vmem[2086] = 8'd116;
vmem[2087] = 8'd105;
vmem[2088] = 8'd115;
vmem[2089] = 8'd32;
vmem[2090] = 8'd117;
vmem[2091] = 8'd114;
vmem[2092] = 8'd110;
vmem[2093] = 8'd97;
vmem[2094] = 8'd44;
vmem[2095] = 8'd32;
vmem[2096] = 8'd105;
vmem[2097] = 8'd100;
vmem[2098] = 8'd32;
vmem[2099] = 8'd109;
vmem[2100] = 8'd97;
vmem[2101] = 8'd108;
vmem[2102] = 8'd101;
vmem[2103] = 8'd115;
vmem[2104] = 8'd117;
vmem[2105] = 8'd97;
vmem[2106] = 8'd100;
vmem[2107] = 8'd97;
vmem[2108] = 8'd32;
vmem[2109] = 8'd100;
vmem[2110] = 8'd117;
vmem[2111] = 8'd105;
vmem[2112] = 8'd32;
vmem[2113] = 8'd100;
vmem[2114] = 8'd105;
vmem[2115] = 8'd99;
vmem[2116] = 8'd116;
vmem[2117] = 8'd117;
vmem[2118] = 8'd109;
vmem[2119] = 8'd32;
vmem[2120] = 8'd118;
vmem[2121] = 8'd105;
vmem[2122] = 8'd116;
vmem[2123] = 8'd97;
vmem[2124] = 8'd101;
vmem[2125] = 8'd46;
vmem[2126] = 8'd32;
vmem[2127] = 8'd80;
vmem[2128] = 8'd114;
vmem[2129] = 8'd111;
vmem[2130] = 8'd105;
vmem[2131] = 8'd110;
vmem[2132] = 8'd32;
vmem[2133] = 8'd114;
vmem[2134] = 8'd117;
vmem[2135] = 8'd116;
vmem[2136] = 8'd114;
vmem[2137] = 8'd117;
vmem[2138] = 8'd109;
vmem[2139] = 8'd32;
vmem[2140] = 8'd114;
vmem[2141] = 8'd105;
vmem[2142] = 8'd115;
vmem[2143] = 8'd117;
vmem[2144] = 8'd115;
vmem[2145] = 8'd32;
vmem[2146] = 8'd97;
vmem[2147] = 8'd99;
vmem[2148] = 8'd32;
vmem[2149] = 8'd102;
vmem[2150] = 8'd101;
vmem[2151] = 8'd108;
vmem[2152] = 8'd105;
vmem[2153] = 8'd115;
vmem[2154] = 8'd32;
vmem[2155] = 8'd111;
vmem[2156] = 8'd114;
vmem[2157] = 8'd110;
vmem[2158] = 8'd97;
vmem[2159] = 8'd114;
vmem[2160] = 8'd101;
vmem[2161] = 8'd32;
vmem[2162] = 8'd102;
vmem[2163] = 8'd114;
vmem[2164] = 8'd105;
vmem[2165] = 8'd110;
vmem[2166] = 8'd103;
vmem[2167] = 8'd105;
vmem[2168] = 8'd108;
vmem[2169] = 8'd108;
vmem[2170] = 8'd97;
vmem[2171] = 8'd46;
vmem[2172] = 8'd32;
vmem[2173] = 8'd68;
vmem[2174] = 8'd111;
vmem[2175] = 8'd110;
vmem[2176] = 8'd101;
vmem[2177] = 8'd99;
vmem[2178] = 8'd32;
vmem[2179] = 8'd101;
vmem[2180] = 8'd108;
vmem[2181] = 8'd101;
vmem[2182] = 8'd109;
vmem[2183] = 8'd101;
vmem[2184] = 8'd110;
vmem[2185] = 8'd116;
vmem[2186] = 8'd117;
vmem[2187] = 8'd109;
vmem[2188] = 8'd32;
vmem[2189] = 8'd108;
vmem[2190] = 8'd101;
vmem[2191] = 8'd99;
vmem[2192] = 8'd116;
vmem[2193] = 8'd117;
vmem[2194] = 8'd115;
vmem[2195] = 8'd32;
vmem[2196] = 8'd113;
vmem[2197] = 8'd117;
vmem[2198] = 8'd97;
vmem[2199] = 8'd109;
vmem[2200] = 8'd44;
vmem[2201] = 8'd32;
vmem[2202] = 8'd105;
vmem[2203] = 8'd110;
vmem[2204] = 8'd32;
vmem[2205] = 8'd112;
vmem[2206] = 8'd101;
vmem[2207] = 8'd108;
vmem[2208] = 8'd108;
vmem[2209] = 8'd101;
vmem[2210] = 8'd110;
vmem[2211] = 8'd116;
vmem[2212] = 8'd101;
vmem[2213] = 8'd115;
vmem[2214] = 8'd113;
vmem[2215] = 8'd117;
vmem[2216] = 8'd101;
vmem[2217] = 8'd32;
vmem[2218] = 8'd108;
vmem[2219] = 8'd101;
vmem[2220] = 8'd111;
vmem[2221] = 8'd32;
vmem[2222] = 8'd117;
vmem[2223] = 8'd108;
vmem[2224] = 8'd116;
vmem[2225] = 8'd114;
vmem[2226] = 8'd105;
vmem[2227] = 8'd99;
vmem[2228] = 8'd105;
vmem[2229] = 8'd101;
vmem[2230] = 8'd115;
vmem[2231] = 8'd32;
vmem[2232] = 8'd97;
vmem[2233] = 8'd116;
vmem[2234] = 8'd46;
vmem[2235] = 8'd32;
vmem[2236] = 8'd73;
vmem[2237] = 8'd110;
vmem[2238] = 8'd32;
vmem[2239] = 8'd116;
vmem[2240] = 8'd105;
vmem[2241] = 8'd110;
vmem[2242] = 8'd99;
vmem[2243] = 8'd105;
vmem[2244] = 8'd100;
vmem[2245] = 8'd117;
vmem[2246] = 8'd110;
vmem[2247] = 8'd116;
vmem[2248] = 8'd32;
vmem[2249] = 8'd116;
vmem[2250] = 8'd105;
vmem[2251] = 8'd110;
vmem[2252] = 8'd99;
vmem[2253] = 8'd105;
vmem[2254] = 8'd100;
vmem[2255] = 8'd117;
vmem[2256] = 8'd110;
vmem[2257] = 8'd116;
vmem[2258] = 8'd32;
vmem[2259] = 8'd101;
vmem[2260] = 8'd102;
vmem[2261] = 8'd102;
vmem[2262] = 8'd105;
vmem[2263] = 8'd99;
vmem[2264] = 8'd105;
vmem[2265] = 8'd116;
vmem[2266] = 8'd117;
vmem[2267] = 8'd114;
vmem[2268] = 8'd46;
vmem[2269] = 8'd32;
vmem[2270] = 8'd68;
vmem[2271] = 8'd111;
vmem[2272] = 8'd110;
vmem[2273] = 8'd101;
vmem[2274] = 8'd99;
vmem[2275] = 8'd32;
vmem[2276] = 8'd97;
vmem[2277] = 8'd99;
vmem[2278] = 8'd99;
vmem[2279] = 8'd117;
vmem[2280] = 8'd109;
vmem[2281] = 8'd115;
vmem[2282] = 8'd97;
vmem[2283] = 8'd110;
vmem[2284] = 8'd44;
vmem[2285] = 8'd32;
vmem[2286] = 8'd102;
vmem[2287] = 8'd101;
vmem[2288] = 8'd108;
vmem[2289] = 8'd105;
vmem[2290] = 8'd115;
vmem[2291] = 8'd32;
vmem[2292] = 8'd108;
vmem[2293] = 8'd97;
vmem[2294] = 8'd99;
vmem[2295] = 8'd105;
vmem[2296] = 8'd110;
vmem[2297] = 8'd105;
vmem[2298] = 8'd97;
vmem[2299] = 8'd32;
vmem[2300] = 8'd100;
vmem[2301] = 8'd105;
vmem[2302] = 8'd103;
vmem[2303] = 8'd110;
vmem[2304] = 8'd105;
vmem[2305] = 8'd115;
vmem[2306] = 8'd115;
vmem[2307] = 8'd105;
vmem[2308] = 8'd109;
vmem[2309] = 8'd32;
vmem[2310] = 8'd116;
vmem[2311] = 8'd101;
vmem[2312] = 8'd109;
vmem[2313] = 8'd112;
vmem[2314] = 8'd111;
vmem[2315] = 8'd114;
vmem[2316] = 8'd44;
vmem[2317] = 8'd32;
vmem[2318] = 8'd115;
vmem[2319] = 8'd101;
vmem[2320] = 8'd109;
vmem[2321] = 8'd32;
vmem[2322] = 8'd113;
vmem[2323] = 8'd117;
vmem[2324] = 8'd97;
vmem[2325] = 8'd109;
vmem[2326] = 8'd32;
vmem[2327] = 8'd109;
vmem[2328] = 8'd97;
vmem[2329] = 8'd108;
vmem[2330] = 8'd101;
vmem[2331] = 8'd115;
vmem[2332] = 8'd117;
vmem[2333] = 8'd97;
vmem[2334] = 8'd100;
vmem[2335] = 8'd97;
vmem[2336] = 8'd32;
vmem[2337] = 8'd108;
vmem[2338] = 8'd111;
vmem[2339] = 8'd114;
vmem[2340] = 8'd101;
vmem[2341] = 8'd109;
vmem[2342] = 8'd44;
vmem[2343] = 8'd32;
vmem[2344] = 8'd117;
vmem[2345] = 8'd108;
vmem[2346] = 8'd116;
vmem[2347] = 8'd114;
vmem[2348] = 8'd105;
vmem[2349] = 8'd99;
vmem[2350] = 8'd101;
vmem[2351] = 8'd115;
vmem[2352] = 8'd32;
vmem[2353] = 8'd115;
vmem[2354] = 8'd117;
vmem[2355] = 8'd115;
vmem[2356] = 8'd99;
vmem[2357] = 8'd105;
vmem[2358] = 8'd112;
vmem[2359] = 8'd105;
vmem[2360] = 8'd116;
vmem[2361] = 8'd32;
vmem[2362] = 8'd110;
vmem[2363] = 8'd117;
vmem[2364] = 8'd110;
vmem[2365] = 8'd99;
vmem[2366] = 8'd32;
vmem[2367] = 8'd101;
vmem[2368] = 8'd120;
vmem[2369] = 8'd32;
vmem[2370] = 8'd101;
vmem[2371] = 8'd116;
vmem[2372] = 8'd32;
vmem[2373] = 8'd101;
vmem[2374] = 8'd120;
vmem[2375] = 8'd46;
vmem[2376] = 8'd32;
vmem[2377] = 8'd86;
vmem[2378] = 8'd101;
vmem[2379] = 8'd115;
vmem[2380] = 8'd116;
vmem[2381] = 8'd105;
vmem[2382] = 8'd98;
vmem[2383] = 8'd117;
vmem[2384] = 8'd108;
vmem[2385] = 8'd117;
vmem[2386] = 8'd109;
vmem[2387] = 8'd32;
vmem[2388] = 8'd97;
vmem[2389] = 8'd116;
vmem[2390] = 8'd32;
vmem[2391] = 8'd116;
vmem[2392] = 8'd101;
vmem[2393] = 8'd109;
vmem[2394] = 8'd112;
vmem[2395] = 8'd111;
vmem[2396] = 8'd114;
vmem[2397] = 8'd32;
vmem[2398] = 8'd101;
vmem[2399] = 8'd120;
vmem[2400] = 8'd44;
vmem[2401] = 8'd32;
vmem[2402] = 8'd115;
vmem[2403] = 8'd105;
vmem[2404] = 8'd116;
vmem[2405] = 8'd32;
vmem[2406] = 8'd97;
vmem[2407] = 8'd109;
vmem[2408] = 8'd101;
vmem[2409] = 8'd116;
vmem[2410] = 8'd32;
vmem[2411] = 8'd109;
vmem[2412] = 8'd97;
vmem[2413] = 8'd108;
vmem[2414] = 8'd101;
vmem[2415] = 8'd115;
vmem[2416] = 8'd117;
vmem[2417] = 8'd97;
vmem[2418] = 8'd100;
vmem[2419] = 8'd97;
vmem[2420] = 8'd32;
vmem[2421] = 8'd106;
vmem[2422] = 8'd117;
vmem[2423] = 8'd115;
vmem[2424] = 8'd116;
vmem[2425] = 8'd111;
vmem[2426] = 8'd46;
vmem[2427] = 8'd32;
vmem[2428] = 8'd73;
vmem[2429] = 8'd110;
vmem[2430] = 8'd116;
vmem[2431] = 8'd101;
vmem[2432] = 8'd103;
vmem[2433] = 8'd101;
vmem[2434] = 8'd114;
vmem[2435] = 8'd32;
vmem[2436] = 8'd97;
vmem[2437] = 8'd108;
vmem[2438] = 8'd105;
vmem[2439] = 8'd113;
vmem[2440] = 8'd117;
vmem[2441] = 8'd101;
vmem[2442] = 8'd116;
vmem[2443] = 8'd32;
vmem[2444] = 8'd111;
vmem[2445] = 8'd114;
vmem[2446] = 8'd110;
vmem[2447] = 8'd97;
vmem[2448] = 8'd114;
vmem[2449] = 8'd101;
vmem[2450] = 8'd32;
vmem[2451] = 8'd109;
vmem[2452] = 8'd97;
vmem[2453] = 8'd117;
vmem[2454] = 8'd114;
vmem[2455] = 8'd105;
vmem[2456] = 8'd115;
vmem[2457] = 8'd32;
vmem[2458] = 8'd105;
vmem[2459] = 8'd110;
vmem[2460] = 8'd32;
vmem[2461] = 8'd118;
vmem[2462] = 8'd101;
vmem[2463] = 8'd110;
vmem[2464] = 8'd101;
vmem[2465] = 8'd110;
vmem[2466] = 8'd97;
vmem[2467] = 8'd116;
vmem[2468] = 8'd105;
vmem[2469] = 8'd115;
vmem[2470] = 8'd46;
vmem[2471] = 8'd32;
vmem[2472] = 8'd85;
vmem[2473] = 8'd116;
vmem[2474] = 8'd32;
vmem[2475] = 8'd101;
vmem[2476] = 8'd117;
vmem[2477] = 8'd32;
vmem[2478] = 8'd110;
vmem[2479] = 8'd101;
vmem[2480] = 8'd113;
vmem[2481] = 8'd117;
vmem[2482] = 8'd101;
vmem[2483] = 8'd32;
vmem[2484] = 8'd101;
vmem[2485] = 8'd117;
vmem[2486] = 8'd32;
vmem[2487] = 8'd109;
vmem[2488] = 8'd97;
vmem[2489] = 8'd103;
vmem[2490] = 8'd110;
vmem[2491] = 8'd97;
vmem[2492] = 8'd32;
vmem[2493] = 8'd115;
vmem[2494] = 8'd101;
vmem[2495] = 8'd109;
vmem[2496] = 8'd112;
vmem[2497] = 8'd101;
vmem[2498] = 8'd114;
vmem[2499] = 8'd32;
vmem[2500] = 8'd102;
vmem[2501] = 8'd97;
vmem[2502] = 8'd99;
vmem[2503] = 8'd105;
vmem[2504] = 8'd108;
vmem[2505] = 8'd105;
vmem[2506] = 8'd115;
vmem[2507] = 8'd105;
vmem[2508] = 8'd115;
vmem[2509] = 8'd46;
vmem[2510] = 8'd32;
vmem[2511] = 8'd83;
vmem[2512] = 8'd117;
vmem[2513] = 8'd115;
vmem[2514] = 8'd112;
vmem[2515] = 8'd101;
vmem[2516] = 8'd110;
vmem[2517] = 8'd100;
vmem[2518] = 8'd105;
vmem[2519] = 8'd115;
vmem[2520] = 8'd115;
vmem[2521] = 8'd101;
vmem[2522] = 8'd32;
vmem[2523] = 8'd109;
vmem[2524] = 8'd101;
vmem[2525] = 8'd116;
vmem[2526] = 8'd117;
vmem[2527] = 8'd115;
vmem[2528] = 8'd32;
vmem[2529] = 8'd111;
vmem[2530] = 8'd100;
vmem[2531] = 8'd105;
vmem[2532] = 8'd111;
vmem[2533] = 8'd44;
vmem[2534] = 8'd32;
vmem[2535] = 8'd101;
vmem[2536] = 8'd102;
vmem[2537] = 8'd102;
vmem[2538] = 8'd105;
vmem[2539] = 8'd99;
vmem[2540] = 8'd105;
vmem[2541] = 8'd116;
vmem[2542] = 8'd117;
vmem[2543] = 8'd114;
vmem[2544] = 8'd32;
vmem[2545] = 8'd110;
vmem[2546] = 8'd101;
vmem[2547] = 8'd99;
vmem[2548] = 8'd32;
vmem[2549] = 8'd102;
vmem[2550] = 8'd114;
vmem[2551] = 8'd105;
vmem[2552] = 8'd110;
vmem[2553] = 8'd103;
vmem[2554] = 8'd105;
vmem[2555] = 8'd108;
vmem[2556] = 8'd108;
vmem[2557] = 8'd97;
vmem[2558] = 8'd32;
vmem[2559] = 8'd105;
vmem[2560] = 8'd110;
vmem[2561] = 8'd44;
vmem[2562] = 8'd32;
vmem[2563] = 8'd115;
vmem[2564] = 8'd111;
vmem[2565] = 8'd108;
vmem[2566] = 8'd108;
vmem[2567] = 8'd105;
vmem[2568] = 8'd99;
vmem[2569] = 8'd105;
vmem[2570] = 8'd116;
vmem[2571] = 8'd117;
vmem[2572] = 8'd100;
vmem[2573] = 8'd105;
vmem[2574] = 8'd110;
vmem[2575] = 8'd32;
vmem[2576] = 8'd115;
vmem[2577] = 8'd97;
vmem[2578] = 8'd103;
vmem[2579] = 8'd105;
vmem[2580] = 8'd116;
vmem[2581] = 8'd116;
vmem[2582] = 8'd105;
vmem[2583] = 8'd115;
vmem[2584] = 8'd32;
vmem[2585] = 8'd116;
vmem[2586] = 8'd117;
vmem[2587] = 8'd114;
vmem[2588] = 8'd112;
vmem[2589] = 8'd105;
vmem[2590] = 8'd115;
vmem[2591] = 8'd46;
vmem[2592] = 8'd32;
vmem[2593] = 8'd73;
vmem[2594] = 8'd110;
vmem[2595] = 8'd32;
vmem[2596] = 8'd112;
vmem[2597] = 8'd101;
vmem[2598] = 8'd108;
vmem[2599] = 8'd108;
vmem[2600] = 8'd101;
vmem[2601] = 8'd110;
vmem[2602] = 8'd116;
vmem[2603] = 8'd101;
vmem[2604] = 8'd115;
vmem[2605] = 8'd113;
vmem[2606] = 8'd117;
vmem[2607] = 8'd101;
vmem[2608] = 8'd32;
vmem[2609] = 8'd108;
vmem[2610] = 8'd117;
vmem[2611] = 8'd99;
vmem[2612] = 8'd116;
vmem[2613] = 8'd117;
vmem[2614] = 8'd115;
vmem[2615] = 8'd32;
vmem[2616] = 8'd99;
vmem[2617] = 8'd111;
vmem[2618] = 8'd110;
vmem[2619] = 8'd115;
vmem[2620] = 8'd101;
vmem[2621] = 8'd113;
vmem[2622] = 8'd117;
vmem[2623] = 8'd97;
vmem[2624] = 8'd116;
vmem[2625] = 8'd46;
vmem[2626] = 8'd32;
vmem[2627] = 8'd67;
vmem[2628] = 8'd114;
vmem[2629] = 8'd97;
vmem[2630] = 8'd115;
vmem[2631] = 8'd32;
vmem[2632] = 8'd115;
vmem[2633] = 8'd111;
vmem[2634] = 8'd100;
vmem[2635] = 8'd97;
vmem[2636] = 8'd108;
vmem[2637] = 8'd101;
vmem[2638] = 8'd115;
vmem[2639] = 8'd32;
vmem[2640] = 8'd116;
vmem[2641] = 8'd111;
vmem[2642] = 8'd114;
vmem[2643] = 8'd116;
vmem[2644] = 8'd111;
vmem[2645] = 8'd114;
vmem[2646] = 8'd32;
vmem[2647] = 8'd117;
vmem[2648] = 8'd108;
vmem[2649] = 8'd116;
vmem[2650] = 8'd114;
vmem[2651] = 8'd105;
vmem[2652] = 8'd99;
vmem[2653] = 8'd105;
vmem[2654] = 8'd101;
vmem[2655] = 8'd115;
vmem[2656] = 8'd44;
vmem[2657] = 8'd32;
vmem[2658] = 8'd102;
vmem[2659] = 8'd114;
vmem[2660] = 8'd105;
vmem[2661] = 8'd110;
vmem[2662] = 8'd103;
vmem[2663] = 8'd105;
vmem[2664] = 8'd108;
vmem[2665] = 8'd108;
vmem[2666] = 8'd97;
vmem[2667] = 8'd32;
vmem[2668] = 8'd110;
vmem[2669] = 8'd117;
vmem[2670] = 8'd108;
vmem[2671] = 8'd108;
vmem[2672] = 8'd97;
vmem[2673] = 8'd32;
vmem[2674] = 8'd97;
vmem[2675] = 8'd99;
vmem[2676] = 8'd44;
vmem[2677] = 8'd32;
vmem[2678] = 8'd98;
vmem[2679] = 8'd105;
vmem[2680] = 8'd98;
vmem[2681] = 8'd101;
vmem[2682] = 8'd110;
vmem[2683] = 8'd100;
vmem[2684] = 8'd117;
vmem[2685] = 8'd109;
vmem[2686] = 8'd32;
vmem[2687] = 8'd100;
vmem[2688] = 8'd117;
vmem[2689] = 8'd105;
vmem[2690] = 8'd46;
vmem[2691] = 8'd32;
vmem[2692] = 8'd67;
vmem[2693] = 8'd117;
vmem[2694] = 8'd114;
vmem[2695] = 8'd97;
vmem[2696] = 8'd98;
vmem[2697] = 8'd105;
vmem[2698] = 8'd116;
vmem[2699] = 8'd117;
vmem[2700] = 8'd114;
vmem[2701] = 8'd32;
vmem[2702] = 8'd101;
vmem[2703] = 8'd103;
vmem[2704] = 8'd101;
vmem[2705] = 8'd115;
vmem[2706] = 8'd116;
vmem[2707] = 8'd97;
vmem[2708] = 8'd115;
vmem[2709] = 8'd32;
vmem[2710] = 8'd109;
vmem[2711] = 8'd97;
vmem[2712] = 8'd120;
vmem[2713] = 8'd105;
vmem[2714] = 8'd109;
vmem[2715] = 8'd117;
vmem[2716] = 8'd115;
vmem[2717] = 8'd32;
vmem[2718] = 8'd108;
vmem[2719] = 8'd101;
vmem[2720] = 8'd111;
vmem[2721] = 8'd32;
vmem[2722] = 8'd112;
vmem[2723] = 8'd111;
vmem[2724] = 8'd114;
vmem[2725] = 8'd116;
vmem[2726] = 8'd116;
vmem[2727] = 8'd105;
vmem[2728] = 8'd116;
vmem[2729] = 8'd111;
vmem[2730] = 8'd114;
vmem[2731] = 8'd32;
vmem[2732] = 8'd109;
vmem[2733] = 8'd111;
vmem[2734] = 8'd108;
vmem[2735] = 8'd101;
vmem[2736] = 8'd115;
vmem[2737] = 8'd116;
vmem[2738] = 8'd105;
vmem[2739] = 8'd101;
vmem[2740] = 8'd46;
vmem[2741] = 8'd32;
vmem[2742] = 8'd86;
vmem[2743] = 8'd101;
vmem[2744] = 8'd115;
vmem[2745] = 8'd116;
vmem[2746] = 8'd105;
vmem[2747] = 8'd98;
vmem[2748] = 8'd117;
vmem[2749] = 8'd108;
vmem[2750] = 8'd117;
vmem[2751] = 8'd109;
vmem[2752] = 8'd32;
vmem[2753] = 8'd101;
vmem[2754] = 8'd115;
vmem[2755] = 8'd116;
vmem[2756] = 8'd32;
vmem[2757] = 8'd97;
vmem[2758] = 8'd110;
vmem[2759] = 8'd116;
vmem[2760] = 8'd101;
vmem[2761] = 8'd44;
vmem[2762] = 8'd32;
vmem[2763] = 8'd99;
vmem[2764] = 8'd111;
vmem[2765] = 8'd110;
vmem[2766] = 8'd100;
vmem[2767] = 8'd105;
vmem[2768] = 8'd109;
vmem[2769] = 8'd101;
vmem[2770] = 8'd110;
vmem[2771] = 8'd116;
vmem[2772] = 8'd117;
vmem[2773] = 8'd109;
vmem[2774] = 8'd32;
vmem[2775] = 8'd97;
vmem[2776] = 8'd32;
vmem[2777] = 8'd108;
vmem[2778] = 8'd101;
vmem[2779] = 8'd99;
vmem[2780] = 8'd116;
vmem[2781] = 8'd117;
vmem[2782] = 8'd115;
vmem[2783] = 8'd32;
vmem[2784] = 8'd113;
vmem[2785] = 8'd117;
vmem[2786] = 8'd105;
vmem[2787] = 8'd115;
vmem[2788] = 8'd44;
vmem[2789] = 8'd32;
vmem[2790] = 8'd108;
vmem[2791] = 8'd97;
vmem[2792] = 8'd111;
vmem[2793] = 8'd114;
vmem[2794] = 8'd101;
vmem[2795] = 8'd101;
vmem[2796] = 8'd116;
vmem[2797] = 8'd32;
vmem[2798] = 8'd116;
vmem[2799] = 8'd101;
vmem[2800] = 8'd109;
vmem[2801] = 8'd112;
vmem[2802] = 8'd117;
vmem[2803] = 8'd115;
vmem[2804] = 8'd32;
vmem[2805] = 8'd108;
vmem[2806] = 8'd101;
vmem[2807] = 8'd111;
vmem[2808] = 8'd46;
vmem[2809] = 8'd32;
vmem[2810] = 8'd76;
vmem[2811] = 8'd111;
vmem[2812] = 8'd114;
vmem[2813] = 8'd101;
vmem[2814] = 8'd109;
vmem[2815] = 8'd32;
vmem[2816] = 8'd105;
vmem[2817] = 8'd112;
vmem[2818] = 8'd115;
vmem[2819] = 8'd117;
vmem[2820] = 8'd109;
vmem[2821] = 8'd32;
vmem[2822] = 8'd100;
vmem[2823] = 8'd111;
vmem[2824] = 8'd108;
vmem[2825] = 8'd111;
vmem[2826] = 8'd114;
vmem[2827] = 8'd32;
vmem[2828] = 8'd115;
vmem[2829] = 8'd105;
vmem[2830] = 8'd116;
vmem[2831] = 8'd32;
vmem[2832] = 8'd97;
vmem[2833] = 8'd109;
vmem[2834] = 8'd101;
vmem[2835] = 8'd116;
vmem[2836] = 8'd44;
vmem[2837] = 8'd32;
vmem[2838] = 8'd99;
vmem[2839] = 8'd111;
vmem[2840] = 8'd110;
vmem[2841] = 8'd115;
vmem[2842] = 8'd101;
vmem[2843] = 8'd99;
vmem[2844] = 8'd116;
vmem[2845] = 8'd101;
vmem[2846] = 8'd116;
vmem[2847] = 8'd117;
vmem[2848] = 8'd114;
vmem[2849] = 8'd32;
vmem[2850] = 8'd97;
vmem[2851] = 8'd100;
vmem[2852] = 8'd105;
vmem[2853] = 8'd112;
vmem[2854] = 8'd105;
vmem[2855] = 8'd115;
vmem[2856] = 8'd99;
vmem[2857] = 8'd105;
vmem[2858] = 8'd110;
vmem[2859] = 8'd103;
vmem[2860] = 8'd32;
vmem[2861] = 8'd101;
vmem[2862] = 8'd108;
vmem[2863] = 8'd105;
vmem[2864] = 8'd116;
vmem[2865] = 8'd46;
vmem[2866] = 8'd32;
vmem[2867] = 8'd80;
vmem[2868] = 8'd101;
vmem[2869] = 8'd108;
vmem[2870] = 8'd108;
vmem[2871] = 8'd101;
vmem[2872] = 8'd110;
vmem[2873] = 8'd116;
vmem[2874] = 8'd101;
vmem[2875] = 8'd115;
vmem[2876] = 8'd113;
vmem[2877] = 8'd117;
vmem[2878] = 8'd101;
vmem[2879] = 8'd32;
vmem[2880] = 8'd118;
vmem[2881] = 8'd111;
vmem[2882] = 8'd108;
vmem[2883] = 8'd117;
vmem[2884] = 8'd116;
vmem[2885] = 8'd112;
vmem[2886] = 8'd97;
vmem[2887] = 8'd116;
vmem[2888] = 8'd32;
vmem[2889] = 8'd115;
vmem[2890] = 8'd111;
vmem[2891] = 8'd108;
vmem[2892] = 8'd108;
vmem[2893] = 8'd105;
vmem[2894] = 8'd99;
vmem[2895] = 8'd105;
vmem[2896] = 8'd116;
vmem[2897] = 8'd117;
vmem[2898] = 8'd100;
vmem[2899] = 8'd105;
vmem[2900] = 8'd110;
vmem[2901] = 8'd32;
vmem[2902] = 8'd111;
vmem[2903] = 8'd100;
vmem[2904] = 8'd105;
vmem[2905] = 8'd111;
vmem[2906] = 8'd32;
vmem[2907] = 8'd105;
vmem[2908] = 8'd100;
vmem[2909] = 8'd32;
vmem[2910] = 8'd115;
vmem[2911] = 8'd101;
vmem[2912] = 8'd109;
vmem[2913] = 8'd112;
vmem[2914] = 8'd101;
vmem[2915] = 8'd114;
vmem[2916] = 8'd46;
vmem[2917] = 8'd32;
vmem[2918] = 8'd73;
vmem[2919] = 8'd110;
vmem[2920] = 8'd116;
vmem[2921] = 8'd101;
vmem[2922] = 8'd114;
vmem[2923] = 8'd100;
vmem[2924] = 8'd117;
vmem[2925] = 8'd109;
vmem[2926] = 8'd32;
vmem[2927] = 8'd101;
vmem[2928] = 8'd116;
vmem[2929] = 8'd32;
vmem[2930] = 8'd109;
vmem[2931] = 8'd97;
vmem[2932] = 8'd108;
vmem[2933] = 8'd101;
vmem[2934] = 8'd115;
vmem[2935] = 8'd117;
vmem[2936] = 8'd97;
vmem[2937] = 8'd100;
vmem[2938] = 8'd97;
vmem[2939] = 8'd32;
vmem[2940] = 8'd102;
vmem[2941] = 8'd97;
vmem[2942] = 8'd109;
vmem[2943] = 8'd101;
vmem[2944] = 8'd115;
vmem[2945] = 8'd32;
vmem[2946] = 8'd97;
vmem[2947] = 8'd99;
vmem[2948] = 8'd32;
vmem[2949] = 8'd97;
vmem[2950] = 8'd110;
vmem[2951] = 8'd116;
vmem[2952] = 8'd101;
vmem[2953] = 8'd32;
vmem[2954] = 8'd105;
vmem[2955] = 8'd112;
vmem[2956] = 8'd115;
vmem[2957] = 8'd117;
vmem[2958] = 8'd109;
vmem[2959] = 8'd32;
vmem[2960] = 8'd112;
vmem[2961] = 8'd114;
vmem[2962] = 8'd105;
vmem[2963] = 8'd109;
vmem[2964] = 8'd105;
vmem[2965] = 8'd115;
vmem[2966] = 8'd32;
vmem[2967] = 8'd105;
vmem[2968] = 8'd110;
vmem[2969] = 8'd32;
vmem[2970] = 8'd102;
vmem[2971] = 8'd97;
vmem[2972] = 8'd117;
vmem[2973] = 8'd99;
vmem[2974] = 8'd105;
vmem[2975] = 8'd98;
vmem[2976] = 8'd117;
vmem[2977] = 8'd115;
vmem[2978] = 8'd46;
vmem[2979] = 8'd32;
vmem[2980] = 8'd65;
vmem[2981] = 8'd108;
vmem[2982] = 8'd105;
vmem[2983] = 8'd113;
vmem[2984] = 8'd117;
vmem[2985] = 8'd97;
vmem[2986] = 8'd109;
vmem[2987] = 8'd32;
vmem[2988] = 8'd114;
vmem[2989] = 8'd117;
vmem[2990] = 8'd116;
vmem[2991] = 8'd114;
vmem[2992] = 8'd117;
vmem[2993] = 8'd109;
vmem[2994] = 8'd32;
vmem[2995] = 8'd99;
vmem[2996] = 8'd111;
vmem[2997] = 8'd110;
vmem[2998] = 8'd115;
vmem[2999] = 8'd101;
vmem[3000] = 8'd113;
vmem[3001] = 8'd117;
vmem[3002] = 8'd97;
vmem[3003] = 8'd116;
vmem[3004] = 8'd32;
vmem[3005] = 8'd118;
vmem[3006] = 8'd101;
vmem[3007] = 8'd108;
vmem[3008] = 8'd105;
vmem[3009] = 8'd116;
vmem[3010] = 8'd32;
vmem[3011] = 8'd113;
vmem[3012] = 8'd117;
vmem[3013] = 8'd105;
vmem[3014] = 8'd115;
vmem[3015] = 8'd32;
vmem[3016] = 8'd101;
vmem[3017] = 8'd108;
vmem[3018] = 8'd101;
vmem[3019] = 8'd105;
vmem[3020] = 8'd102;
vmem[3021] = 8'd101;
vmem[3022] = 8'd110;
vmem[3023] = 8'd100;
vmem[3024] = 8'd46;
vmem[3025] = 8'd32;
vmem[3026] = 8'd67;
vmem[3027] = 8'd117;
vmem[3028] = 8'd114;
vmem[3029] = 8'd97;
vmem[3030] = 8'd98;
vmem[3031] = 8'd105;
vmem[3032] = 8'd116;
vmem[3033] = 8'd117;
vmem[3034] = 8'd114;
vmem[3035] = 8'd32;
vmem[3036] = 8'd97;
vmem[3037] = 8'd108;
vmem[3038] = 8'd105;
vmem[3039] = 8'd113;
vmem[3040] = 8'd117;
vmem[3041] = 8'd101;
vmem[3042] = 8'd116;
vmem[3043] = 8'd32;
vmem[3044] = 8'd108;
vmem[3045] = 8'd117;
vmem[3046] = 8'd99;
vmem[3047] = 8'd116;
vmem[3048] = 8'd117;
vmem[3049] = 8'd115;
vmem[3050] = 8'd32;
vmem[3051] = 8'd116;
vmem[3052] = 8'd101;
vmem[3053] = 8'd108;
vmem[3054] = 8'd108;
vmem[3055] = 8'd117;
vmem[3056] = 8'd115;
vmem[3057] = 8'd32;
vmem[3058] = 8'd97;
vmem[3059] = 8'd116;
vmem[3060] = 8'd32;
vmem[3061] = 8'd112;
vmem[3062] = 8'd111;
vmem[3063] = 8'd115;
vmem[3064] = 8'd117;
vmem[3065] = 8'd101;
vmem[3066] = 8'd114;
vmem[3067] = 8'd101;
vmem[3068] = 8'd46;
vmem[3069] = 8'd32;
vmem[3070] = 8'd78;
vmem[3071] = 8'd97;
vmem[3072] = 8'd109;
vmem[3073] = 8'd32;
vmem[3074] = 8'd103;
vmem[3075] = 8'd114;
vmem[3076] = 8'd97;
vmem[3077] = 8'd118;
vmem[3078] = 8'd105;
vmem[3079] = 8'd100;
vmem[3080] = 8'd97;
vmem[3081] = 8'd32;
vmem[3082] = 8'd108;
vmem[3083] = 8'd105;
vmem[3084] = 8'd98;
vmem[3085] = 8'd101;
vmem[3086] = 8'd114;
vmem[3087] = 8'd111;
vmem[3088] = 8'd32;
vmem[3089] = 8'd97;
vmem[3090] = 8'd99;
vmem[3091] = 8'd32;
vmem[3092] = 8'd108;
vmem[3093] = 8'd117;
vmem[3094] = 8'd99;
vmem[3095] = 8'd116;
vmem[3096] = 8'd117;
vmem[3097] = 8'd115;
vmem[3098] = 8'd32;
vmem[3099] = 8'd105;
vmem[3100] = 8'd110;
vmem[3101] = 8'd116;
vmem[3102] = 8'd101;
vmem[3103] = 8'd114;
vmem[3104] = 8'd100;
vmem[3105] = 8'd117;
vmem[3106] = 8'd109;
vmem[3107] = 8'd46;
vmem[3108] = 8'd32;
vmem[3109] = 8'd83;
vmem[3110] = 8'd101;
vmem[3111] = 8'd100;
vmem[3112] = 8'd32;
vmem[3113] = 8'd117;
vmem[3114] = 8'd108;
vmem[3115] = 8'd116;
vmem[3116] = 8'd114;
vmem[3117] = 8'd105;
vmem[3118] = 8'd99;
vmem[3119] = 8'd101;
vmem[3120] = 8'd115;
vmem[3121] = 8'd32;
vmem[3122] = 8'd109;
vmem[3123] = 8'd105;
vmem[3124] = 8'd32;
vmem[3125] = 8'd110;
vmem[3126] = 8'd111;
vmem[3127] = 8'd110;
vmem[3128] = 8'd32;
vmem[3129] = 8'd118;
vmem[3130] = 8'd101;
vmem[3131] = 8'd108;
vmem[3132] = 8'd105;
vmem[3133] = 8'd116;
vmem[3134] = 8'd32;
vmem[3135] = 8'd101;
vmem[3136] = 8'd117;
vmem[3137] = 8'd105;
vmem[3138] = 8'd115;
vmem[3139] = 8'd109;
vmem[3140] = 8'd111;
vmem[3141] = 8'd100;
vmem[3142] = 8'd32;
vmem[3143] = 8'd112;
vmem[3144] = 8'd101;
vmem[3145] = 8'd108;
vmem[3146] = 8'd108;
vmem[3147] = 8'd101;
vmem[3148] = 8'd110;
vmem[3149] = 8'd116;
vmem[3150] = 8'd101;
vmem[3151] = 8'd115;
vmem[3152] = 8'd113;
vmem[3153] = 8'd117;
vmem[3154] = 8'd101;
vmem[3155] = 8'd46;
vmem[3156] = 8'd32;
vmem[3157] = 8'd67;
vmem[3158] = 8'd108;
vmem[3159] = 8'd97;
vmem[3160] = 8'd115;
vmem[3161] = 8'd115;
vmem[3162] = 8'd32;
vmem[3163] = 8'd97;
vmem[3164] = 8'd112;
vmem[3165] = 8'd116;
vmem[3166] = 8'd101;
vmem[3167] = 8'd110;
vmem[3168] = 8'd116;
vmem[3169] = 8'd32;
vmem[3170] = 8'd116;
vmem[3171] = 8'd97;
vmem[3172] = 8'd99;
vmem[3173] = 8'd105;
vmem[3174] = 8'd116;
vmem[3175] = 8'd105;
vmem[3176] = 8'd32;
vmem[3177] = 8'd115;
vmem[3178] = 8'd111;
vmem[3179] = 8'd99;
vmem[3180] = 8'd105;
vmem[3181] = 8'd111;
vmem[3182] = 8'd115;
vmem[3183] = 8'd113;
vmem[3184] = 8'd117;
vmem[3185] = 8'd32;
vmem[3186] = 8'd97;
vmem[3187] = 8'd100;
vmem[3188] = 8'd32;
vmem[3189] = 8'd108;
vmem[3190] = 8'd105;
vmem[3191] = 8'd116;
vmem[3192] = 8'd111;
vmem[3193] = 8'd114;
vmem[3194] = 8'd97;
vmem[3195] = 8'd32;
vmem[3196] = 8'd116;
vmem[3197] = 8'd111;
vmem[3198] = 8'd114;
vmem[3199] = 8'd113;
vmem[3200] = 8'd117;
vmem[3201] = 8'd101;
vmem[3202] = 8'd110;
vmem[3203] = 8'd116;
vmem[3204] = 8'd32;
vmem[3205] = 8'd112;
vmem[3206] = 8'd101;
vmem[3207] = 8'd114;
vmem[3208] = 8'd32;
vmem[3209] = 8'd99;
vmem[3210] = 8'd111;
vmem[3211] = 8'd110;
vmem[3212] = 8'd117;
vmem[3213] = 8'd98;
vmem[3214] = 8'd105;
vmem[3215] = 8'd97;
vmem[3216] = 8'd32;
vmem[3217] = 8'd110;
vmem[3218] = 8'd111;
vmem[3219] = 8'd115;
vmem[3220] = 8'd116;
vmem[3221] = 8'd114;
vmem[3222] = 8'd97;
vmem[3223] = 8'd44;
vmem[3224] = 8'd32;
vmem[3225] = 8'd112;
vmem[3226] = 8'd101;
vmem[3227] = 8'd114;
vmem[3228] = 8'd32;
vmem[3229] = 8'd105;
vmem[3230] = 8'd110;
vmem[3231] = 8'd99;
vmem[3232] = 8'd101;
vmem[3233] = 8'd112;
vmem[3234] = 8'd116;
vmem[3235] = 8'd111;
vmem[3236] = 8'd115;
vmem[3237] = 8'd32;
vmem[3238] = 8'd104;
vmem[3239] = 8'd105;
vmem[3240] = 8'd109;
vmem[3241] = 8'd101;
vmem[3242] = 8'd110;
vmem[3243] = 8'd97;
vmem[3244] = 8'd101;
vmem[3245] = 8'd111;
vmem[3246] = 8'd115;
vmem[3247] = 8'd46;
vmem[3248] = 8'd32;
vmem[3249] = 8'd83;
vmem[3250] = 8'd117;
vmem[3251] = 8'd115;
vmem[3252] = 8'd112;
vmem[3253] = 8'd101;
vmem[3254] = 8'd110;
vmem[3255] = 8'd100;
vmem[3256] = 8'd105;
vmem[3257] = 8'd115;
vmem[3258] = 8'd115;
vmem[3259] = 8'd101;
vmem[3260] = 8'd32;
vmem[3261] = 8'd97;
vmem[3262] = 8'd108;
vmem[3263] = 8'd105;
vmem[3264] = 8'd113;
vmem[3265] = 8'd117;
vmem[3266] = 8'd97;
vmem[3267] = 8'd109;
vmem[3268] = 8'd32;
vmem[3269] = 8'd101;
vmem[3270] = 8'd108;
vmem[3271] = 8'd101;
vmem[3272] = 8'd105;
vmem[3273] = 8'd102;
vmem[3274] = 8'd101;
vmem[3275] = 8'd110;
vmem[3276] = 8'd100;
vmem[3277] = 8'd32;
vmem[3278] = 8'd102;
vmem[3279] = 8'd101;
vmem[3280] = 8'd114;
vmem[3281] = 8'd109;
vmem[3282] = 8'd101;
vmem[3283] = 8'd110;
vmem[3284] = 8'd116;
vmem[3285] = 8'd117;
vmem[3286] = 8'd109;
vmem[3287] = 8'd46;
vmem[3288] = 8'd32;
vmem[3289] = 8'd73;
vmem[3290] = 8'd110;
vmem[3291] = 8'd32;
vmem[3292] = 8'd115;
vmem[3293] = 8'd117;
vmem[3294] = 8'd115;
vmem[3295] = 8'd99;
vmem[3296] = 8'd105;
vmem[3297] = 8'd112;
vmem[3298] = 8'd105;
vmem[3299] = 8'd116;
vmem[3300] = 8'd32;
vmem[3301] = 8'd100;
vmem[3302] = 8'd105;
vmem[3303] = 8'd103;
vmem[3304] = 8'd110;
vmem[3305] = 8'd105;
vmem[3306] = 8'd115;
vmem[3307] = 8'd115;
vmem[3308] = 8'd105;
vmem[3309] = 8'd109;
vmem[3310] = 8'd32;
vmem[3311] = 8'd105;
vmem[3312] = 8'd110;
vmem[3313] = 8'd116;
vmem[3314] = 8'd101;
vmem[3315] = 8'd114;
vmem[3316] = 8'd100;
vmem[3317] = 8'd117;
vmem[3318] = 8'd109;
vmem[3319] = 8'd46;
vmem[3320] = 8'd32;
vmem[3321] = 8'd67;
vmem[3322] = 8'd114;
vmem[3323] = 8'd97;
vmem[3324] = 8'd115;
vmem[3325] = 8'd32;
vmem[3326] = 8'd100;
vmem[3327] = 8'd105;
vmem[3328] = 8'd103;
vmem[3329] = 8'd110;
vmem[3330] = 8'd105;
vmem[3331] = 8'd115;
vmem[3332] = 8'd115;
vmem[3333] = 8'd105;
vmem[3334] = 8'd109;
vmem[3335] = 8'd32;
vmem[3336] = 8'd111;
vmem[3337] = 8'd114;
vmem[3338] = 8'd99;
vmem[3339] = 8'd105;
vmem[3340] = 8'd32;
vmem[3341] = 8'd101;
vmem[3342] = 8'd103;
vmem[3343] = 8'd101;
vmem[3344] = 8'd116;
vmem[3345] = 8'd32;
vmem[3346] = 8'd116;
vmem[3347] = 8'd114;
vmem[3348] = 8'd105;
vmem[3349] = 8'd115;
vmem[3350] = 8'd116;
vmem[3351] = 8'd105;
vmem[3352] = 8'd113;
vmem[3353] = 8'd117;
vmem[3354] = 8'd101;
vmem[3355] = 8'd32;
vmem[3356] = 8'd116;
vmem[3357] = 8'd101;
vmem[3358] = 8'd109;
vmem[3359] = 8'd112;
vmem[3360] = 8'd111;
vmem[3361] = 8'd114;
vmem[3362] = 8'd46;
vmem[3363] = 8'd32;
vmem[3364] = 8'd83;
vmem[3365] = 8'd117;
vmem[3366] = 8'd115;
vmem[3367] = 8'd112;
vmem[3368] = 8'd101;
vmem[3369] = 8'd110;
vmem[3370] = 8'd100;
vmem[3371] = 8'd105;
vmem[3372] = 8'd115;
vmem[3373] = 8'd115;
vmem[3374] = 8'd101;
vmem[3375] = 8'd32;
vmem[3376] = 8'd97;
vmem[3377] = 8'd99;
vmem[3378] = 8'd32;
vmem[3379] = 8'd116;
vmem[3380] = 8'd101;
vmem[3381] = 8'd108;
vmem[3382] = 8'd108;
vmem[3383] = 8'd117;
vmem[3384] = 8'd115;
vmem[3385] = 8'd32;
vmem[3386] = 8'd115;
vmem[3387] = 8'd111;
vmem[3388] = 8'd108;
vmem[3389] = 8'd108;
vmem[3390] = 8'd105;
vmem[3391] = 8'd99;
vmem[3392] = 8'd105;
vmem[3393] = 8'd116;
vmem[3394] = 8'd117;
vmem[3395] = 8'd100;
vmem[3396] = 8'd105;
vmem[3397] = 8'd110;
vmem[3398] = 8'd44;
vmem[3399] = 8'd32;
vmem[3400] = 8'd118;
vmem[3401] = 8'd105;
vmem[3402] = 8'd118;
vmem[3403] = 8'd101;
vmem[3404] = 8'd114;
vmem[3405] = 8'd114;
vmem[3406] = 8'd97;
vmem[3407] = 8'd32;
vmem[3408] = 8'd100;
vmem[3409] = 8'd105;
vmem[3410] = 8'd97;
vmem[3411] = 8'd109;
vmem[3412] = 8'd32;
vmem[3413] = 8'd105;
vmem[3414] = 8'd100;
vmem[3415] = 8'd44;
vmem[3416] = 8'd32;
vmem[3417] = 8'd112;
vmem[3418] = 8'd101;
vmem[3419] = 8'd108;
vmem[3420] = 8'd108;
vmem[3421] = 8'd101;
vmem[3422] = 8'd110;
vmem[3423] = 8'd116;
vmem[3424] = 8'd101;
vmem[3425] = 8'd115;
vmem[3426] = 8'd113;
vmem[3427] = 8'd117;
vmem[3428] = 8'd101;
vmem[3429] = 8'd32;
vmem[3430] = 8'd109;
vmem[3431] = 8'd97;
vmem[3432] = 8'd103;
vmem[3433] = 8'd110;
vmem[3434] = 8'd97;
vmem[3435] = 8'd46;
vmem[3436] = 8'd32;
vmem[3437] = 8'd86;
vmem[3438] = 8'd105;
vmem[3439] = 8'd118;
vmem[3440] = 8'd97;
vmem[3441] = 8'd109;
vmem[3442] = 8'd117;
vmem[3443] = 8'd115;
vmem[3444] = 8'd32;
vmem[3445] = 8'd112;
vmem[3446] = 8'd111;
vmem[3447] = 8'd114;
vmem[3448] = 8'd116;
vmem[3449] = 8'd116;
vmem[3450] = 8'd105;
vmem[3451] = 8'd116;
vmem[3452] = 8'd111;
vmem[3453] = 8'd114;
vmem[3454] = 8'd32;
vmem[3455] = 8'd108;
vmem[3456] = 8'd101;
vmem[3457] = 8'd111;
vmem[3458] = 8'd32;
vmem[3459] = 8'd100;
vmem[3460] = 8'd105;
vmem[3461] = 8'd97;
vmem[3462] = 8'd109;
vmem[3463] = 8'd44;
vmem[3464] = 8'd32;
vmem[3465] = 8'd101;
vmem[3466] = 8'd117;
vmem[3467] = 8'd32;
vmem[3468] = 8'd117;
vmem[3469] = 8'd108;
vmem[3470] = 8'd116;
vmem[3471] = 8'd114;
vmem[3472] = 8'd105;
vmem[3473] = 8'd99;
vmem[3474] = 8'd105;
vmem[3475] = 8'd101;
vmem[3476] = 8'd115;
vmem[3477] = 8'd32;
vmem[3478] = 8'd116;
vmem[3479] = 8'd101;
vmem[3480] = 8'd108;
vmem[3481] = 8'd108;
vmem[3482] = 8'd117;
vmem[3483] = 8'd115;
vmem[3484] = 8'd32;
vmem[3485] = 8'd118;
vmem[3486] = 8'd111;
vmem[3487] = 8'd108;
vmem[3488] = 8'd117;
vmem[3489] = 8'd116;
vmem[3490] = 8'd112;
vmem[3491] = 8'd97;
vmem[3492] = 8'd116;
vmem[3493] = 8'd32;
vmem[3494] = 8'd97;
vmem[3495] = 8'd46;
vmem[3496] = 8'd32;
vmem[3497] = 8'd67;
vmem[3498] = 8'd114;
vmem[3499] = 8'd97;
vmem[3500] = 8'd115;
vmem[3501] = 8'd32;
vmem[3502] = 8'd99;
vmem[3503] = 8'd111;
vmem[3504] = 8'd110;
vmem[3505] = 8'd115;
vmem[3506] = 8'd101;
vmem[3507] = 8'd113;
vmem[3508] = 8'd117;
vmem[3509] = 8'd97;
vmem[3510] = 8'd116;
vmem[3511] = 8'd32;
vmem[3512] = 8'd110;
vmem[3513] = 8'd105;
vmem[3514] = 8'd115;
vmem[3515] = 8'd108;
vmem[3516] = 8'd32;
vmem[3517] = 8'd118;
vmem[3518] = 8'd105;
vmem[3519] = 8'd116;
vmem[3520] = 8'd97;
vmem[3521] = 8'd101;
vmem[3522] = 8'd32;
vmem[3523] = 8'd117;
vmem[3524] = 8'd114;
vmem[3525] = 8'd110;
vmem[3526] = 8'd97;
vmem[3527] = 8'd32;
vmem[3528] = 8'd99;
vmem[3529] = 8'd117;
vmem[3530] = 8'd114;
vmem[3531] = 8'd115;
vmem[3532] = 8'd117;
vmem[3533] = 8'd115;
vmem[3534] = 8'd32;
vmem[3535] = 8'd101;
vmem[3536] = 8'd108;
vmem[3537] = 8'd101;
vmem[3538] = 8'd105;
vmem[3539] = 8'd102;
vmem[3540] = 8'd101;
vmem[3541] = 8'd110;
vmem[3542] = 8'd100;
vmem[3543] = 8'd46;
vmem[3544] = 8'd32;
vmem[3545] = 8'd67;
vmem[3546] = 8'd114;
vmem[3547] = 8'd97;
vmem[3548] = 8'd115;
vmem[3549] = 8'd32;
vmem[3550] = 8'd117;
vmem[3551] = 8'd108;
vmem[3552] = 8'd116;
vmem[3553] = 8'd114;
vmem[3554] = 8'd105;
vmem[3555] = 8'd99;
vmem[3556] = 8'd105;
vmem[3557] = 8'd101;
vmem[3558] = 8'd115;
vmem[3559] = 8'd32;
vmem[3560] = 8'd97;
vmem[3561] = 8'd117;
vmem[3562] = 8'd103;
vmem[3563] = 8'd117;
vmem[3564] = 8'd101;
vmem[3565] = 8'd32;
vmem[3566] = 8'd97;
vmem[3567] = 8'd116;
vmem[3568] = 8'd32;
vmem[3569] = 8'd100;
vmem[3570] = 8'd111;
vmem[3571] = 8'd108;
vmem[3572] = 8'd111;
vmem[3573] = 8'd114;
vmem[3574] = 8'd32;
vmem[3575] = 8'd102;
vmem[3576] = 8'd97;
vmem[3577] = 8'd99;
vmem[3578] = 8'd105;
vmem[3579] = 8'd108;
vmem[3580] = 8'd105;
vmem[3581] = 8'd115;
vmem[3582] = 8'd105;
vmem[3583] = 8'd115;
vmem[3584] = 8'd32;
vmem[3585] = 8'd118;
vmem[3586] = 8'd105;
vmem[3587] = 8'd118;
vmem[3588] = 8'd101;
vmem[3589] = 8'd114;
vmem[3590] = 8'd114;
vmem[3591] = 8'd97;
vmem[3592] = 8'd46;
vmem[3593] = 8'd32;
vmem[3594] = 8'd70;
vmem[3595] = 8'd117;
vmem[3596] = 8'd115;
vmem[3597] = 8'd99;
vmem[3598] = 8'd101;
vmem[3599] = 8'd32;
vmem[3600] = 8'd109;
vmem[3601] = 8'd105;
vmem[3602] = 8'd32;
vmem[3603] = 8'd116;
vmem[3604] = 8'd101;
vmem[3605] = 8'd108;
vmem[3606] = 8'd108;
vmem[3607] = 8'd117;
vmem[3608] = 8'd115;
vmem[3609] = 8'd44;
vmem[3610] = 8'd32;
vmem[3611] = 8'd118;
vmem[3612] = 8'd111;
vmem[3613] = 8'd108;
vmem[3614] = 8'd117;
vmem[3615] = 8'd116;
vmem[3616] = 8'd112;
vmem[3617] = 8'd97;
vmem[3618] = 8'd116;
vmem[3619] = 8'd32;
vmem[3620] = 8'd102;
vmem[3621] = 8'd101;
vmem[3622] = 8'd114;
vmem[3623] = 8'd109;
vmem[3624] = 8'd101;
vmem[3625] = 8'd110;
vmem[3626] = 8'd116;
vmem[3627] = 8'd117;
vmem[3628] = 8'd109;
vmem[3629] = 8'd32;
vmem[3630] = 8'd97;
vmem[3631] = 8'd114;
vmem[3632] = 8'd99;
vmem[3633] = 8'd117;
vmem[3634] = 8'd32;
vmem[3635] = 8'd108;
vmem[3636] = 8'd111;
vmem[3637] = 8'd98;
vmem[3638] = 8'd111;
vmem[3639] = 8'd114;
vmem[3640] = 8'd116;
vmem[3641] = 8'd105;
vmem[3642] = 8'd115;
vmem[3643] = 8'd44;
vmem[3644] = 8'd32;
vmem[3645] = 8'd104;
vmem[3646] = 8'd101;
vmem[3647] = 8'd110;
vmem[3648] = 8'd100;
vmem[3649] = 8'd114;
vmem[3650] = 8'd101;
vmem[3651] = 8'd114;
vmem[3652] = 8'd105;
vmem[3653] = 8'd116;
vmem[3654] = 8'd32;
vmem[3655] = 8'd112;
vmem[3656] = 8'd111;
vmem[3657] = 8'd114;
vmem[3658] = 8'd116;
vmem[3659] = 8'd97;
vmem[3660] = 8'd32;
vmem[3661] = 8'd110;
vmem[3662] = 8'd101;
vmem[3663] = 8'd113;
vmem[3664] = 8'd117;
vmem[3665] = 8'd101;
vmem[3666] = 8'd46;
vmem[3667] = 8'd32;
vmem[3668] = 8'd80;
vmem[3669] = 8'd114;
vmem[3670] = 8'd111;
vmem[3671] = 8'd105;
vmem[3672] = 8'd110;
vmem[3673] = 8'd32;
vmem[3674] = 8'd117;
vmem[3675] = 8'd116;
vmem[3676] = 8'd32;
vmem[3677] = 8'd109;
vmem[3678] = 8'd97;
vmem[3679] = 8'd115;
vmem[3680] = 8'd115;
vmem[3681] = 8'd97;
vmem[3682] = 8'd32;
vmem[3683] = 8'd118;
vmem[3684] = 8'd105;
vmem[3685] = 8'd116;
vmem[3686] = 8'd97;
vmem[3687] = 8'd101;
vmem[3688] = 8'd32;
vmem[3689] = 8'd115;
vmem[3690] = 8'd101;
vmem[3691] = 8'd109;
vmem[3692] = 8'd32;
vmem[3693] = 8'd112;
vmem[3694] = 8'd108;
vmem[3695] = 8'd97;
vmem[3696] = 8'd99;
vmem[3697] = 8'd101;
vmem[3698] = 8'd114;
vmem[3699] = 8'd97;
vmem[3700] = 8'd116;
vmem[3701] = 8'd32;
vmem[3702] = 8'd99;
vmem[3703] = 8'd111;
vmem[3704] = 8'd109;
vmem[3705] = 8'd109;
vmem[3706] = 8'd111;
vmem[3707] = 8'd100;
vmem[3708] = 8'd111;
vmem[3709] = 8'd32;
vmem[3710] = 8'd115;
vmem[3711] = 8'd101;
vmem[3712] = 8'd100;
vmem[3713] = 8'd32;
vmem[3714] = 8'd101;
vmem[3715] = 8'd116;
vmem[3716] = 8'd32;
vmem[3717] = 8'd108;
vmem[3718] = 8'd101;
vmem[3719] = 8'd111;
vmem[3720] = 8'd46;
vmem[3721] = 8'd32;
vmem[3722] = 8'd78;
vmem[3723] = 8'd117;
vmem[3724] = 8'd108;
vmem[3725] = 8'd108;
vmem[3726] = 8'd97;
vmem[3727] = 8'd109;
vmem[3728] = 8'd32;
vmem[3729] = 8'd98;
vmem[3730] = 8'd105;
vmem[3731] = 8'd98;
vmem[3732] = 8'd101;
vmem[3733] = 8'd110;
vmem[3734] = 8'd100;
vmem[3735] = 8'd117;
vmem[3736] = 8'd109;
vmem[3737] = 8'd32;
vmem[3738] = 8'd97;
vmem[3739] = 8'd117;
vmem[3740] = 8'd103;
vmem[3741] = 8'd117;
vmem[3742] = 8'd101;
vmem[3743] = 8'd32;
vmem[3744] = 8'd101;
vmem[3745] = 8'd116;
vmem[3746] = 8'd32;
vmem[3747] = 8'd108;
vmem[3748] = 8'd101;
vmem[3749] = 8'd99;
vmem[3750] = 8'd116;
vmem[3751] = 8'd117;
vmem[3752] = 8'd115;
vmem[3753] = 8'd32;
vmem[3754] = 8'd112;
vmem[3755] = 8'd111;
vmem[3756] = 8'd114;
vmem[3757] = 8'd116;
vmem[3758] = 8'd116;
vmem[3759] = 8'd105;
vmem[3760] = 8'd116;
vmem[3761] = 8'd111;
vmem[3762] = 8'd114;
vmem[3763] = 8'd32;
vmem[3764] = 8'd117;
vmem[3765] = 8'd108;
vmem[3766] = 8'd116;
vmem[3767] = 8'd114;
vmem[3768] = 8'd105;
vmem[3769] = 8'd99;
vmem[3770] = 8'd101;
vmem[3771] = 8'd115;
vmem[3772] = 8'd46;
vmem[3773] = 8'd32;
vmem[3774] = 8'd78;
vmem[3775] = 8'd117;
vmem[3776] = 8'd110;
vmem[3777] = 8'd99;
vmem[3778] = 8'd32;
vmem[3779] = 8'd116;
vmem[3780] = 8'd101;
vmem[3781] = 8'd109;
vmem[3782] = 8'd112;
vmem[3783] = 8'd111;
vmem[3784] = 8'd114;
vmem[3785] = 8'd32;
vmem[3786] = 8'd109;
vmem[3787] = 8'd101;
vmem[3788] = 8'd116;
vmem[3789] = 8'd117;
vmem[3790] = 8'd115;
vmem[3791] = 8'd32;
vmem[3792] = 8'd118;
vmem[3793] = 8'd101;
vmem[3794] = 8'd108;
vmem[3795] = 8'd32;
vmem[3796] = 8'd111;
vmem[3797] = 8'd100;
vmem[3798] = 8'd105;
vmem[3799] = 8'd111;
vmem[3800] = 8'd32;
vmem[3801] = 8'd99;
vmem[3802] = 8'd111;
vmem[3803] = 8'd110;
vmem[3804] = 8'd103;
vmem[3805] = 8'd117;
vmem[3806] = 8'd101;
vmem[3807] = 8'd32;
vmem[3808] = 8'd116;
vmem[3809] = 8'd114;
vmem[3810] = 8'd105;
vmem[3811] = 8'd115;
vmem[3812] = 8'd116;
vmem[3813] = 8'd105;
vmem[3814] = 8'd113;
vmem[3815] = 8'd117;
vmem[3816] = 8'd101;
vmem[3817] = 8'd46;
vmem[3818] = 8'd32;
vmem[3819] = 8'd78;
vmem[3820] = 8'd97;
vmem[3821] = 8'd109;
vmem[3822] = 8'd32;
vmem[3823] = 8'd108;
vmem[3824] = 8'd105;
vmem[3825] = 8'd103;
vmem[3826] = 8'd117;
vmem[3827] = 8'd108;
vmem[3828] = 8'd97;
vmem[3829] = 8'd32;
vmem[3830] = 8'd111;
vmem[3831] = 8'd100;
vmem[3832] = 8'd105;
vmem[3833] = 8'd111;
vmem[3834] = 8'd44;
vmem[3835] = 8'd32;
vmem[3836] = 8'd102;
vmem[3837] = 8'd97;
vmem[3838] = 8'd99;
vmem[3839] = 8'd105;
vmem[3840] = 8'd108;
vmem[3841] = 8'd105;
vmem[3842] = 8'd115;
vmem[3843] = 8'd105;
vmem[3844] = 8'd115;
vmem[3845] = 8'd32;
vmem[3846] = 8'd118;
vmem[3847] = 8'd101;
vmem[3848] = 8'd108;
vmem[3849] = 8'd32;
vmem[3850] = 8'd108;
vmem[3851] = 8'd97;
vmem[3852] = 8'd111;
vmem[3853] = 8'd114;
vmem[3854] = 8'd101;
vmem[3855] = 8'd101;
vmem[3856] = 8'd116;
vmem[3857] = 8'd32;
vmem[3858] = 8'd101;
vmem[3859] = 8'd103;
vmem[3860] = 8'd101;
vmem[3861] = 8'd116;
vmem[3862] = 8'd44;
vmem[3863] = 8'd32;
vmem[3864] = 8'd99;
vmem[3865] = 8'd111;
vmem[3866] = 8'd110;
vmem[3867] = 8'd118;
vmem[3868] = 8'd97;
vmem[3869] = 8'd108;
vmem[3870] = 8'd108;
vmem[3871] = 8'd105;
vmem[3872] = 8'd115;
vmem[3873] = 8'd32;
vmem[3874] = 8'd110;
vmem[3875] = 8'd111;
vmem[3876] = 8'd110;
vmem[3877] = 8'd32;
vmem[3878] = 8'd108;
vmem[3879] = 8'd105;
vmem[3880] = 8'd98;
vmem[3881] = 8'd101;
vmem[3882] = 8'd114;
vmem[3883] = 8'd111;
vmem[3884] = 8'd46;
vmem[3885] = 8'd32;
vmem[3886] = 8'd80;
vmem[3887] = 8'd101;
vmem[3888] = 8'd108;
vmem[3889] = 8'd108;
vmem[3890] = 8'd101;
vmem[3891] = 8'd110;
vmem[3892] = 8'd116;
vmem[3893] = 8'd101;
vmem[3894] = 8'd115;
vmem[3895] = 8'd113;
vmem[3896] = 8'd117;
vmem[3897] = 8'd101;
vmem[3898] = 8'd32;
vmem[3899] = 8'd105;
vmem[3900] = 8'd110;
vmem[3901] = 8'd32;
vmem[3902] = 8'd108;
vmem[3903] = 8'd111;
vmem[3904] = 8'd114;
vmem[3905] = 8'd101;
vmem[3906] = 8'd109;
vmem[3907] = 8'd32;
vmem[3908] = 8'd115;
vmem[3909] = 8'd105;
vmem[3910] = 8'd116;
vmem[3911] = 8'd32;
vmem[3912] = 8'd97;
vmem[3913] = 8'd109;
vmem[3914] = 8'd101;
vmem[3915] = 8'd116;
vmem[3916] = 8'd32;
vmem[3917] = 8'd118;
vmem[3918] = 8'd101;
vmem[3919] = 8'd108;
vmem[3920] = 8'd105;
vmem[3921] = 8'd116;
vmem[3922] = 8'd32;
vmem[3923] = 8'd109;
vmem[3924] = 8'd111;
vmem[3925] = 8'd108;
vmem[3926] = 8'd101;
vmem[3927] = 8'd115;
vmem[3928] = 8'd116;
vmem[3929] = 8'd105;
vmem[3930] = 8'd101;
vmem[3931] = 8'd32;
vmem[3932] = 8'd99;
vmem[3933] = 8'd111;
vmem[3934] = 8'd110;
vmem[3935] = 8'd103;
vmem[3936] = 8'd117;
vmem[3937] = 8'd101;
vmem[3938] = 8'd32;
vmem[3939] = 8'd97;
vmem[3940] = 8'd32;
vmem[3941] = 8'd115;
vmem[3942] = 8'd105;
vmem[3943] = 8'd116;
vmem[3944] = 8'd32;
vmem[3945] = 8'd97;
vmem[3946] = 8'd109;
vmem[3947] = 8'd101;
vmem[3948] = 8'd116;
vmem[3949] = 8'd32;
vmem[3950] = 8'd113;
vmem[3951] = 8'd117;
vmem[3952] = 8'd97;
vmem[3953] = 8'd109;
vmem[3954] = 8'd46;
vmem[3955] = 8'd32;
vmem[3956] = 8'd83;
vmem[3957] = 8'd101;
vmem[3958] = 8'd100;
vmem[3959] = 8'd32;
vmem[3960] = 8'd115;
vmem[3961] = 8'd101;
vmem[3962] = 8'd100;
vmem[3963] = 8'd32;
vmem[3964] = 8'd100;
vmem[3965] = 8'd105;
vmem[3966] = 8'd99;
vmem[3967] = 8'd116;
vmem[3968] = 8'd117;
vmem[3969] = 8'd109;
vmem[3970] = 8'd32;
vmem[3971] = 8'd110;
vmem[3972] = 8'd101;
vmem[3973] = 8'd113;
vmem[3974] = 8'd117;
vmem[3975] = 8'd101;
vmem[3976] = 8'd44;
vmem[3977] = 8'd32;
vmem[3978] = 8'd97;
vmem[3979] = 8'd117;
vmem[3980] = 8'd99;
vmem[3981] = 8'd116;
vmem[3982] = 8'd111;
vmem[3983] = 8'd114;
vmem[3984] = 8'd32;
vmem[3985] = 8'd117;
vmem[3986] = 8'd108;
vmem[3987] = 8'd108;
vmem[3988] = 8'd97;
vmem[3989] = 8'd109;
vmem[3990] = 8'd99;
vmem[3991] = 8'd111;
vmem[3992] = 8'd114;
vmem[3993] = 8'd112;
vmem[3994] = 8'd101;
vmem[3995] = 8'd114;
vmem[3996] = 8'd32;
vmem[3997] = 8'd114;
vmem[3998] = 8'd105;
vmem[3999] = 8'd115;
vmem[4000] = 8'd117;
vmem[4001] = 8'd115;
vmem[4002] = 8'd46;
vmem[4003] = 8'd32;
vmem[4004] = 8'd65;
vmem[4005] = 8'd101;
vmem[4006] = 8'd110;
vmem[4007] = 8'd101;
vmem[4008] = 8'd97;
vmem[4009] = 8'd110;
vmem[4010] = 8'd32;
vmem[4011] = 8'd105;
vmem[4012] = 8'd110;
vmem[4013] = 8'd32;
vmem[4014] = 8'd102;
vmem[4015] = 8'd101;
vmem[4016] = 8'd108;
vmem[4017] = 8'd105;
vmem[4018] = 8'd115;
vmem[4019] = 8'd32;
vmem[4020] = 8'd113;
vmem[4021] = 8'd117;
vmem[4022] = 8'd105;
vmem[4023] = 8'd115;
vmem[4024] = 8'd32;
vmem[4025] = 8'd109;
vmem[4026] = 8'd97;
vmem[4027] = 8'd115;
vmem[4028] = 8'd115;
vmem[4029] = 8'd97;
vmem[4030] = 8'd32;
vmem[4031] = 8'd108;
vmem[4032] = 8'd117;
vmem[4033] = 8'd99;
vmem[4034] = 8'd116;
vmem[4035] = 8'd117;
vmem[4036] = 8'd115;
vmem[4037] = 8'd32;
vmem[4038] = 8'd99;
vmem[4039] = 8'd111;
vmem[4040] = 8'd110;
vmem[4041] = 8'd100;
vmem[4042] = 8'd105;
vmem[4043] = 8'd109;
vmem[4044] = 8'd101;
vmem[4045] = 8'd110;
vmem[4046] = 8'd116;
vmem[4047] = 8'd117;
vmem[4048] = 8'd109;
vmem[4049] = 8'd32;
vmem[4050] = 8'd97;
vmem[4051] = 8'd32;
vmem[4052] = 8'd118;
vmem[4053] = 8'd101;
vmem[4054] = 8'd108;
vmem[4055] = 8'd32;
vmem[4056] = 8'd101;
vmem[4057] = 8'd120;
vmem[4058] = 8'd46;
vmem[4059] = 8'd32;
vmem[4060] = 8'd68;
vmem[4061] = 8'd111;
vmem[4062] = 8'd110;
vmem[4063] = 8'd101;
vmem[4064] = 8'd99;
vmem[4065] = 8'd32;
vmem[4066] = 8'd97;
vmem[4067] = 8'd116;
vmem[4068] = 8'd32;
vmem[4069] = 8'd102;
vmem[4070] = 8'd101;
vmem[4071] = 8'd117;
vmem[4072] = 8'd103;
vmem[4073] = 8'd105;
vmem[4074] = 8'd97;
vmem[4075] = 8'd116;
vmem[4076] = 8'd32;
vmem[4077] = 8'd108;
vmem[4078] = 8'd105;
vmem[4079] = 8'd98;
vmem[4080] = 8'd101;
vmem[4081] = 8'd114;
vmem[4082] = 8'd111;
vmem[4083] = 8'd44;
vmem[4084] = 8'd32;
vmem[4085] = 8'd117;
vmem[4086] = 8'd116;
vmem[4087] = 8'd32;
vmem[4088] = 8'd99;
vmem[4089] = 8'd111;
vmem[4090] = 8'd110;
vmem[4091] = 8'd103;
vmem[4092] = 8'd117;
vmem[4093] = 8'd101;
vmem[4094] = 8'd32;
vmem[4095] = 8'd101;
vmem[4096] = 8'd114;
vmem[4097] = 8'd97;
vmem[4098] = 8'd116;
vmem[4099] = 8'd46;
vmem[4100] = 8'd32;
vmem[4101] = 8'd78;
vmem[4102] = 8'd97;
vmem[4103] = 8'd109;
vmem[4104] = 8'd32;
vmem[4105] = 8'd118;
vmem[4106] = 8'd117;
vmem[4107] = 8'd108;
vmem[4108] = 8'd112;
vmem[4109] = 8'd117;
vmem[4110] = 8'd116;
vmem[4111] = 8'd97;
vmem[4112] = 8'd116;
vmem[4113] = 8'd101;
vmem[4114] = 8'd32;
vmem[4115] = 8'd109;
vmem[4116] = 8'd97;
vmem[4117] = 8'd103;
vmem[4118] = 8'd110;
vmem[4119] = 8'd97;
vmem[4120] = 8'd32;
vmem[4121] = 8'd118;
vmem[4122] = 8'd105;
vmem[4123] = 8'd116;
vmem[4124] = 8'd97;
vmem[4125] = 8'd101;
vmem[4126] = 8'd32;
vmem[4127] = 8'd108;
vmem[4128] = 8'd105;
vmem[4129] = 8'd98;
vmem[4130] = 8'd101;
vmem[4131] = 8'd114;
vmem[4132] = 8'd111;
vmem[4133] = 8'd32;
vmem[4134] = 8'd102;
vmem[4135] = 8'd105;
vmem[4136] = 8'd110;
vmem[4137] = 8'd105;
vmem[4138] = 8'd98;
vmem[4139] = 8'd117;
vmem[4140] = 8'd115;
vmem[4141] = 8'd32;
vmem[4142] = 8'd102;
vmem[4143] = 8'd105;
vmem[4144] = 8'd110;
vmem[4145] = 8'd105;
vmem[4146] = 8'd98;
vmem[4147] = 8'd117;
vmem[4148] = 8'd115;
vmem[4149] = 8'd46;
vmem[4150] = 8'd32;
vmem[4151] = 8'd65;
vmem[4152] = 8'd108;
vmem[4153] = 8'd105;
vmem[4154] = 8'd113;
vmem[4155] = 8'd117;
vmem[4156] = 8'd97;
vmem[4157] = 8'd109;
vmem[4158] = 8'd32;
vmem[4159] = 8'd115;
vmem[4160] = 8'd111;
vmem[4161] = 8'd108;
vmem[4162] = 8'd108;
vmem[4163] = 8'd105;
vmem[4164] = 8'd99;
vmem[4165] = 8'd105;
vmem[4166] = 8'd116;
vmem[4167] = 8'd117;
vmem[4168] = 8'd100;
vmem[4169] = 8'd105;
vmem[4170] = 8'd110;
vmem[4171] = 8'd32;
vmem[4172] = 8'd100;
vmem[4173] = 8'd105;
vmem[4174] = 8'd97;
vmem[4175] = 8'd109;
vmem[4176] = 8'd32;
vmem[4177] = 8'd97;
vmem[4178] = 8'd116;
vmem[4179] = 8'd32;
vmem[4180] = 8'd109;
vmem[4181] = 8'd97;
vmem[4182] = 8'd116;
vmem[4183] = 8'd116;
vmem[4184] = 8'd105;
vmem[4185] = 8'd115;
vmem[4186] = 8'd32;
vmem[4187] = 8'd105;
vmem[4188] = 8'd97;
vmem[4189] = 8'd99;
vmem[4190] = 8'd117;
vmem[4191] = 8'd108;
vmem[4192] = 8'd105;
vmem[4193] = 8'd115;
vmem[4194] = 8'd46;
vmem[4195] = 8'd32;
vmem[4196] = 8'd69;
vmem[4197] = 8'd116;
vmem[4198] = 8'd105;
vmem[4199] = 8'd97;
vmem[4200] = 8'd109;
vmem[4201] = 8'd32;
vmem[4202] = 8'd97;
vmem[4203] = 8'd116;
vmem[4204] = 8'd32;
vmem[4205] = 8'd110;
vmem[4206] = 8'd101;
vmem[4207] = 8'd113;
vmem[4208] = 8'd117;
vmem[4209] = 8'd101;
vmem[4210] = 8'd32;
vmem[4211] = 8'd101;
vmem[4212] = 8'd102;
vmem[4213] = 8'd102;
vmem[4214] = 8'd105;
vmem[4215] = 8'd99;
vmem[4216] = 8'd105;
vmem[4217] = 8'd116;
vmem[4218] = 8'd117;
vmem[4219] = 8'd114;
vmem[4220] = 8'd44;
vmem[4221] = 8'd32;
vmem[4222] = 8'd109;
vmem[4223] = 8'd97;
vmem[4224] = 8'd108;
vmem[4225] = 8'd101;
vmem[4226] = 8'd115;
vmem[4227] = 8'd117;
vmem[4228] = 8'd97;
vmem[4229] = 8'd100;
vmem[4230] = 8'd97;
vmem[4231] = 8'd32;
vmem[4232] = 8'd109;
vmem[4233] = 8'd97;
vmem[4234] = 8'd117;
vmem[4235] = 8'd114;
vmem[4236] = 8'd105;
vmem[4237] = 8'd115;
vmem[4238] = 8'd32;
vmem[4239] = 8'd97;
vmem[4240] = 8'd44;
vmem[4241] = 8'd32;
vmem[4242] = 8'd115;
vmem[4243] = 8'd99;
vmem[4244] = 8'd101;
vmem[4245] = 8'd108;
vmem[4246] = 8'd101;
vmem[4247] = 8'd114;
vmem[4248] = 8'd105;
vmem[4249] = 8'd115;
vmem[4250] = 8'd113;
vmem[4251] = 8'd117;
vmem[4252] = 8'd101;
vmem[4253] = 8'd32;
vmem[4254] = 8'd101;
vmem[4255] = 8'd108;
vmem[4256] = 8'd105;
vmem[4257] = 8'd116;
vmem[4258] = 8'd46;
vmem[4259] = 8'd32;
vmem[4260] = 8'd69;
vmem[4261] = 8'd116;
vmem[4262] = 8'd105;
vmem[4263] = 8'd97;
vmem[4264] = 8'd109;
vmem[4265] = 8'd32;
vmem[4266] = 8'd110;
vmem[4267] = 8'd117;
vmem[4268] = 8'd108;
vmem[4269] = 8'd108;
vmem[4270] = 8'd97;
vmem[4271] = 8'd32;
vmem[4272] = 8'd100;
vmem[4273] = 8'd105;
vmem[4274] = 8'd97;
vmem[4275] = 8'd109;
vmem[4276] = 8'd44;
vmem[4277] = 8'd32;
vmem[4278] = 8'd115;
vmem[4279] = 8'd111;
vmem[4280] = 8'd100;
vmem[4281] = 8'd97;
vmem[4282] = 8'd108;
vmem[4283] = 8'd101;
vmem[4284] = 8'd115;
vmem[4285] = 8'd32;
vmem[4286] = 8'd97;
vmem[4287] = 8'd32;
vmem[4288] = 8'd109;
vmem[4289] = 8'd97;
vmem[4290] = 8'd117;
vmem[4291] = 8'd114;
vmem[4292] = 8'd105;
vmem[4293] = 8'd115;
vmem[4294] = 8'd32;
vmem[4295] = 8'd115;
vmem[4296] = 8'd111;
vmem[4297] = 8'd108;
vmem[4298] = 8'd108;
vmem[4299] = 8'd105;
vmem[4300] = 8'd99;
vmem[4301] = 8'd105;
vmem[4302] = 8'd116;
vmem[4303] = 8'd117;
vmem[4304] = 8'd100;
vmem[4305] = 8'd105;
vmem[4306] = 8'd110;
vmem[4307] = 8'd44;
vmem[4308] = 8'd32;
vmem[4309] = 8'd104;
vmem[4310] = 8'd101;
vmem[4311] = 8'd110;
vmem[4312] = 8'd100;
vmem[4313] = 8'd114;
vmem[4314] = 8'd101;
vmem[4315] = 8'd114;
vmem[4316] = 8'd105;
vmem[4317] = 8'd116;
vmem[4318] = 8'd32;
vmem[4319] = 8'd114;
vmem[4320] = 8'd104;
vmem[4321] = 8'd111;
vmem[4322] = 8'd110;
vmem[4323] = 8'd99;
vmem[4324] = 8'd117;
vmem[4325] = 8'd115;
vmem[4326] = 8'd32;
vmem[4327] = 8'd100;
vmem[4328] = 8'd105;
vmem[4329] = 8'd97;
vmem[4330] = 8'd109;
vmem[4331] = 8'd46;
vmem[4332] = 8'd32;
vmem[4333] = 8'd68;
vmem[4334] = 8'd111;
vmem[4335] = 8'd110;
vmem[4336] = 8'd101;
vmem[4337] = 8'd99;
vmem[4338] = 8'd32;
vmem[4339] = 8'd108;
vmem[4340] = 8'd117;
vmem[4341] = 8'd99;
vmem[4342] = 8'd116;
vmem[4343] = 8'd117;
vmem[4344] = 8'd115;
vmem[4345] = 8'd32;
vmem[4346] = 8'd110;
vmem[4347] = 8'd105;
vmem[4348] = 8'd98;
vmem[4349] = 8'd104;
vmem[4350] = 8'd32;
vmem[4351] = 8'd97;
vmem[4352] = 8'd99;
vmem[4353] = 8'd32;
vmem[4354] = 8'd117;
vmem[4355] = 8'd114;
vmem[4356] = 8'd110;
vmem[4357] = 8'd97;
vmem[4358] = 8'd32;
vmem[4359] = 8'd115;
vmem[4360] = 8'd117;
vmem[4361] = 8'd115;
vmem[4362] = 8'd99;
vmem[4363] = 8'd105;
vmem[4364] = 8'd112;
vmem[4365] = 8'd105;
vmem[4366] = 8'd116;
vmem[4367] = 8'd44;
vmem[4368] = 8'd32;
vmem[4369] = 8'd105;
vmem[4370] = 8'd100;
vmem[4371] = 8'd32;
vmem[4372] = 8'd109;
vmem[4373] = 8'd97;
vmem[4374] = 8'd108;
vmem[4375] = 8'd101;
vmem[4376] = 8'd115;
vmem[4377] = 8'd117;
vmem[4378] = 8'd97;
vmem[4379] = 8'd100;
vmem[4380] = 8'd97;
vmem[4381] = 8'd32;
vmem[4382] = 8'd101;
vmem[4383] = 8'd114;
vmem[4384] = 8'd97;
vmem[4385] = 8'd116;
vmem[4386] = 8'd32;
vmem[4387] = 8'd101;
vmem[4388] = 8'd108;
vmem[4389] = 8'd101;
vmem[4390] = 8'd109;
vmem[4391] = 8'd101;
vmem[4392] = 8'd110;
vmem[4393] = 8'd116;
vmem[4394] = 8'd117;
vmem[4395] = 8'd109;
vmem[4396] = 8'd46;
vmem[4397] = 8'd32;
vmem[4398] = 8'd65;
vmem[4399] = 8'd108;
vmem[4400] = 8'd105;
vmem[4401] = 8'd113;
vmem[4402] = 8'd117;
vmem[4403] = 8'd97;
vmem[4404] = 8'd109;
vmem[4405] = 8'd32;
vmem[4406] = 8'd112;
vmem[4407] = 8'd111;
vmem[4408] = 8'd115;
vmem[4409] = 8'd117;
vmem[4410] = 8'd101;
vmem[4411] = 8'd114;
vmem[4412] = 8'd101;
vmem[4413] = 8'd32;
vmem[4414] = 8'd109;
vmem[4415] = 8'd97;
vmem[4416] = 8'd117;
vmem[4417] = 8'd114;
vmem[4418] = 8'd105;
vmem[4419] = 8'd115;
vmem[4420] = 8'd32;
vmem[4421] = 8'd108;
vmem[4422] = 8'd111;
vmem[4423] = 8'd98;
vmem[4424] = 8'd111;
vmem[4425] = 8'd114;
vmem[4426] = 8'd116;
vmem[4427] = 8'd105;
vmem[4428] = 8'd115;
vmem[4429] = 8'd32;
vmem[4430] = 8'd102;
vmem[4431] = 8'd101;
vmem[4432] = 8'd117;
vmem[4433] = 8'd103;
vmem[4434] = 8'd105;
vmem[4435] = 8'd97;
vmem[4436] = 8'd116;
vmem[4437] = 8'd32;
vmem[4438] = 8'd109;
vmem[4439] = 8'd97;
vmem[4440] = 8'd116;
vmem[4441] = 8'd116;
vmem[4442] = 8'd105;
vmem[4443] = 8'd115;
vmem[4444] = 8'd46;
vmem[4445] = 8'd32;
vmem[4446] = 8'd85;
vmem[4447] = 8'd116;
vmem[4448] = 8'd32;
vmem[4449] = 8'd110;
vmem[4450] = 8'd101;
vmem[4451] = 8'd99;
vmem[4452] = 8'd32;
vmem[4453] = 8'd109;
vmem[4454] = 8'd97;
vmem[4455] = 8'd103;
vmem[4456] = 8'd110;
vmem[4457] = 8'd97;
vmem[4458] = 8'd32;
vmem[4459] = 8'd118;
vmem[4460] = 8'd101;
vmem[4461] = 8'd108;
vmem[4462] = 8'd105;
vmem[4463] = 8'd116;
vmem[4464] = 8'd46;
vmem[4465] = 8'd32;
vmem[4466] = 8'd83;
vmem[4467] = 8'd117;
vmem[4468] = 8'd115;
vmem[4469] = 8'd112;
vmem[4470] = 8'd101;
vmem[4471] = 8'd110;
vmem[4472] = 8'd100;
vmem[4473] = 8'd105;
vmem[4474] = 8'd115;
vmem[4475] = 8'd115;
vmem[4476] = 8'd101;
vmem[4477] = 8'd32;
vmem[4478] = 8'd105;
vmem[4479] = 8'd100;
vmem[4480] = 8'd32;
vmem[4481] = 8'd109;
vmem[4482] = 8'd97;
vmem[4483] = 8'd103;
vmem[4484] = 8'd110;
vmem[4485] = 8'd97;
vmem[4486] = 8'd32;
vmem[4487] = 8'd101;
vmem[4488] = 8'd103;
vmem[4489] = 8'd101;
vmem[4490] = 8'd116;
vmem[4491] = 8'd32;
vmem[4492] = 8'd100;
vmem[4493] = 8'd117;
vmem[4494] = 8'd105;
vmem[4495] = 8'd32;
vmem[4496] = 8'd105;
vmem[4497] = 8'd109;
vmem[4498] = 8'd112;
vmem[4499] = 8'd101;
vmem[4500] = 8'd114;
vmem[4501] = 8'd100;
vmem[4502] = 8'd105;
vmem[4503] = 8'd101;
vmem[4504] = 8'd116;
vmem[4505] = 8'd32;
vmem[4506] = 8'd99;
vmem[4507] = 8'd111;
vmem[4508] = 8'd110;
vmem[4509] = 8'd103;
vmem[4510] = 8'd117;
vmem[4511] = 8'd101;
vmem[4512] = 8'd32;
vmem[4513] = 8'd118;
vmem[4514] = 8'd105;
vmem[4515] = 8'd116;
vmem[4516] = 8'd97;
vmem[4517] = 8'd101;
vmem[4518] = 8'd32;
vmem[4519] = 8'd97;
vmem[4520] = 8'd116;
vmem[4521] = 8'd32;
vmem[4522] = 8'd108;
vmem[4523] = 8'd111;
vmem[4524] = 8'd114;
vmem[4525] = 8'd101;
vmem[4526] = 8'd109;
vmem[4527] = 8'd46;
vmem[4528] = 8'd32;
vmem[4529] = 8'd73;
vmem[4530] = 8'd110;
vmem[4531] = 8'd32;
vmem[4532] = 8'd110;
vmem[4533] = 8'd111;
vmem[4534] = 8'd110;
vmem[4535] = 8'd32;
vmem[4536] = 8'd99;
vmem[4537] = 8'd111;
vmem[4538] = 8'd109;
vmem[4539] = 8'd109;
vmem[4540] = 8'd111;
vmem[4541] = 8'd100;
vmem[4542] = 8'd111;
vmem[4543] = 8'd32;
vmem[4544] = 8'd100;
vmem[4545] = 8'd111;
vmem[4546] = 8'd108;
vmem[4547] = 8'd111;
vmem[4548] = 8'd114;
vmem[4549] = 8'd44;
vmem[4550] = 8'd32;
vmem[4551] = 8'd113;
vmem[4552] = 8'd117;
vmem[4553] = 8'd105;
vmem[4554] = 8'd115;
vmem[4555] = 8'd32;
vmem[4556] = 8'd108;
vmem[4557] = 8'd97;
vmem[4558] = 8'd99;
vmem[4559] = 8'd105;
vmem[4560] = 8'd110;
vmem[4561] = 8'd105;
vmem[4562] = 8'd97;
vmem[4563] = 8'd32;
vmem[4564] = 8'd102;
vmem[4565] = 8'd101;
vmem[4566] = 8'd108;
vmem[4567] = 8'd105;
vmem[4568] = 8'd115;
vmem[4569] = 8'd46;
vmem[4570] = 8'd32;
vmem[4571] = 8'd78;
vmem[4572] = 8'd117;
vmem[4573] = 8'd108;
vmem[4574] = 8'd108;
vmem[4575] = 8'd97;
vmem[4576] = 8'd109;
vmem[4577] = 8'd32;
vmem[4578] = 8'd118;
vmem[4579] = 8'd97;
vmem[4580] = 8'd114;
vmem[4581] = 8'd105;
vmem[4582] = 8'd117;
vmem[4583] = 8'd115;
vmem[4584] = 8'd32;
vmem[4585] = 8'd118;
vmem[4586] = 8'd101;
vmem[4587] = 8'd108;
vmem[4588] = 8'd105;
vmem[4589] = 8'd116;
vmem[4590] = 8'd32;
vmem[4591] = 8'd115;
vmem[4592] = 8'd105;
vmem[4593] = 8'd116;
vmem[4594] = 8'd32;
vmem[4595] = 8'd97;
vmem[4596] = 8'd109;
vmem[4597] = 8'd101;
vmem[4598] = 8'd116;
vmem[4599] = 8'd32;
vmem[4600] = 8'd110;
vmem[4601] = 8'd105;
vmem[4602] = 8'd115;
vmem[4603] = 8'd108;
vmem[4604] = 8'd32;
vmem[4605] = 8'd104;
vmem[4606] = 8'd101;
vmem[4607] = 8'd110;
vmem[4608] = 8'd100;
vmem[4609] = 8'd114;
vmem[4610] = 8'd101;
vmem[4611] = 8'd114;
vmem[4612] = 8'd105;
vmem[4613] = 8'd116;
vmem[4614] = 8'd32;
vmem[4615] = 8'd112;
vmem[4616] = 8'd108;
vmem[4617] = 8'd97;
vmem[4618] = 8'd99;
vmem[4619] = 8'd101;
vmem[4620] = 8'd114;
vmem[4621] = 8'd97;
vmem[4622] = 8'd116;
vmem[4623] = 8'd46;
vmem[4624] = 8'd32;
vmem[4625] = 8'd77;
vmem[4626] = 8'd111;
vmem[4627] = 8'd114;
vmem[4628] = 8'd98;
vmem[4629] = 8'd105;
vmem[4630] = 8'd32;
vmem[4631] = 8'd116;
vmem[4632] = 8'd101;
vmem[4633] = 8'd109;
vmem[4634] = 8'd112;
vmem[4635] = 8'd117;
vmem[4636] = 8'd115;
vmem[4637] = 8'd32;
vmem[4638] = 8'd115;
vmem[4639] = 8'd97;
vmem[4640] = 8'd112;
vmem[4641] = 8'd105;
vmem[4642] = 8'd101;
vmem[4643] = 8'd110;
vmem[4644] = 8'd32;
vmem[4645] = 8'd100;
vmem[4646] = 8'd117;
vmem[4647] = 8'd105;
vmem[4648] = 8'd44;
vmem[4649] = 8'd32;
vmem[4650] = 8'd110;
vmem[4651] = 8'd111;
vmem[4652] = 8'd110;
vmem[4653] = 8'd32;
vmem[4654] = 8'd118;
vmem[4655] = 8'd97;
vmem[4656] = 8'd114;
vmem[4657] = 8'd105;
vmem[4658] = 8'd117;
vmem[4659] = 8'd115;
vmem[4660] = 8'd32;
vmem[4661] = 8'd100;
vmem[4662] = 8'd105;
vmem[4663] = 8'd97;
vmem[4664] = 8'd109;
vmem[4665] = 8'd32;
vmem[4666] = 8'd116;
vmem[4667] = 8'd101;
vmem[4668] = 8'd109;
vmem[4669] = 8'd112;
vmem[4670] = 8'd117;
vmem[4671] = 8'd115;
vmem[4672] = 8'd32;
vmem[4673] = 8'd97;
vmem[4674] = 8'd99;
vmem[4675] = 8'd46;
vmem[4676] = 8'd32;
vmem[4677] = 8'd80;
vmem[4678] = 8'd101;
vmem[4679] = 8'd108;
vmem[4680] = 8'd108;
vmem[4681] = 8'd101;
vmem[4682] = 8'd110;
vmem[4683] = 8'd116;
vmem[4684] = 8'd101;
vmem[4685] = 8'd115;
vmem[4686] = 8'd113;
vmem[4687] = 8'd117;
vmem[4688] = 8'd101;
vmem[4689] = 8'd32;
vmem[4690] = 8'd110;
vmem[4691] = 8'd117;
vmem[4692] = 8'd108;
vmem[4693] = 8'd108;
vmem[4694] = 8'd97;
vmem[4695] = 8'd32;
vmem[4696] = 8'd109;
vmem[4697] = 8'd105;
vmem[4698] = 8'd44;
vmem[4699] = 8'd32;
vmem[4700] = 8'd112;
vmem[4701] = 8'd101;
vmem[4702] = 8'd108;
vmem[4703] = 8'd108;
vmem[4704] = 8'd101;
vmem[4705] = 8'd110;
vmem[4706] = 8'd116;
vmem[4707] = 8'd101;
vmem[4708] = 8'd115;
vmem[4709] = 8'd113;
vmem[4710] = 8'd117;
vmem[4711] = 8'd101;
vmem[4712] = 8'd32;
vmem[4713] = 8'd118;
vmem[4714] = 8'd101;
vmem[4715] = 8'd108;
vmem[4716] = 8'd32;
vmem[4717] = 8'd108;
vmem[4718] = 8'd105;
vmem[4719] = 8'd98;
vmem[4720] = 8'd101;
vmem[4721] = 8'd114;
vmem[4722] = 8'd111;
vmem[4723] = 8'd32;
vmem[4724] = 8'd97;
vmem[4725] = 8'd99;
vmem[4726] = 8'd44;
vmem[4727] = 8'd32;
vmem[4728] = 8'd97;
vmem[4729] = 8'd108;
vmem[4730] = 8'd105;
vmem[4731] = 8'd113;
vmem[4732] = 8'd117;
vmem[4733] = 8'd101;
vmem[4734] = 8'd116;
vmem[4735] = 8'd32;
vmem[4736] = 8'd100;
vmem[4737] = 8'd105;
vmem[4738] = 8'd99;
vmem[4739] = 8'd116;
vmem[4740] = 8'd117;
vmem[4741] = 8'd109;
vmem[4742] = 8'd32;
vmem[4743] = 8'd109;
vmem[4744] = 8'd105;
vmem[4745] = 8'd46;
vmem[4746] = 8'd32;
vmem[4747] = 8'd85;
vmem[4748] = 8'd116;
vmem[4749] = 8'd32;
vmem[4750] = 8'd105;
vmem[4751] = 8'd110;
vmem[4752] = 8'd32;
vmem[4753] = 8'd110;
vmem[4754] = 8'd117;
vmem[4755] = 8'd108;
vmem[4756] = 8'd108;
vmem[4757] = 8'd97;
vmem[4758] = 8'd32;
vmem[4759] = 8'd97;
vmem[4760] = 8'd110;
vmem[4761] = 8'd116;
vmem[4762] = 8'd101;
vmem[4763] = 8'd46;
vmem[4764] = 8'd32;
vmem[4765] = 8'd80;
vmem[4766] = 8'd104;
vmem[4767] = 8'd97;
vmem[4768] = 8'd115;
vmem[4769] = 8'd101;
vmem[4770] = 8'd108;
vmem[4771] = 8'd108;
vmem[4772] = 8'd117;
vmem[4773] = 8'd115;
vmem[4774] = 8'd32;
vmem[4775] = 8'd101;
vmem[4776] = 8'd116;
vmem[4777] = 8'd32;
vmem[4778] = 8'd112;
vmem[4779] = 8'd114;
vmem[4780] = 8'd101;
vmem[4781] = 8'd116;
vmem[4782] = 8'd105;
vmem[4783] = 8'd117;
vmem[4784] = 8'd109;
vmem[4785] = 8'd32;
vmem[4786] = 8'd112;
vmem[4787] = 8'd117;
vmem[4788] = 8'd114;
vmem[4789] = 8'd117;
vmem[4790] = 8'd115;
vmem[4791] = 8'd44;
vmem[4792] = 8'd32;
vmem[4793] = 8'd97;
vmem[4794] = 8'd116;
vmem[4795] = 8'd32;
vmem[4796] = 8'd108;
vmem[4797] = 8'd117;
vmem[4798] = 8'd99;
vmem[4799] = 8'd116;
vmem[4800] = 8'd117;
vmem[4801] = 8'd115;
vmem[4802] = 8'd32;
vmem[4803] = 8'd114;
vmem[4804] = 8'd105;
vmem[4805] = 8'd115;
vmem[4806] = 8'd117;
vmem[4807] = 8'd115;
vmem[4808] = 8'd46;
vmem[4809] = 8'd32;
vmem[4810] = 8'd68;
vmem[4811] = 8'd117;
vmem[4812] = 8'd105;
vmem[4813] = 8'd115;
vmem[4814] = 8'd32;
vmem[4815] = 8'd118;
vmem[4816] = 8'd101;
vmem[4817] = 8'd108;
vmem[4818] = 8'd105;
vmem[4819] = 8'd116;
vmem[4820] = 8'd32;
vmem[4821] = 8'd111;
vmem[4822] = 8'd114;
vmem[4823] = 8'd99;
vmem[4824] = 8'd105;
vmem[4825] = 8'd44;
vmem[4826] = 8'd32;
vmem[4827] = 8'd99;
vmem[4828] = 8'd111;
vmem[4829] = 8'd110;
vmem[4830] = 8'd103;
vmem[4831] = 8'd117;
vmem[4832] = 8'd101;
vmem[4833] = 8'd32;
vmem[4834] = 8'd117;
vmem[4835] = 8'd116;
vmem[4836] = 8'd32;
vmem[4837] = 8'd108;
vmem[4838] = 8'd97;
vmem[4839] = 8'd99;
vmem[4840] = 8'd105;
vmem[4841] = 8'd110;
vmem[4842] = 8'd105;
vmem[4843] = 8'd97;
vmem[4844] = 8'd32;
vmem[4845] = 8'd101;
vmem[4846] = 8'd116;
vmem[4847] = 8'd44;
vmem[4848] = 8'd32;
vmem[4849] = 8'd118;
vmem[4850] = 8'd101;
vmem[4851] = 8'd115;
vmem[4852] = 8'd116;
vmem[4853] = 8'd105;
vmem[4854] = 8'd98;
vmem[4855] = 8'd117;
vmem[4856] = 8'd108;
vmem[4857] = 8'd117;
vmem[4858] = 8'd109;
vmem[4859] = 8'd32;
vmem[4860] = 8'd101;
vmem[4861] = 8'd116;
vmem[4862] = 8'd32;
vmem[4863] = 8'd109;
vmem[4864] = 8'd97;
vmem[4865] = 8'd117;
vmem[4866] = 8'd114;
vmem[4867] = 8'd105;
vmem[4868] = 8'd115;
vmem[4869] = 8'd46;
vmem[4870] = 8'd32;
vmem[4871] = 8'd80;
vmem[4872] = 8'd114;
vmem[4873] = 8'd97;
vmem[4874] = 8'd101;
vmem[4875] = 8'd115;
vmem[4876] = 8'd101;
vmem[4877] = 8'd110;
vmem[4878] = 8'd116;
vmem[4879] = 8'd32;
vmem[4880] = 8'd97;
vmem[4881] = 8'd117;
vmem[4882] = 8'd99;
vmem[4883] = 8'd116;
vmem[4884] = 8'd111;
vmem[4885] = 8'd114;
vmem[4886] = 8'd32;
vmem[4887] = 8'd118;
vmem[4888] = 8'd101;
vmem[4889] = 8'd108;
vmem[4890] = 8'd105;
vmem[4891] = 8'd116;
vmem[4892] = 8'd32;
vmem[4893] = 8'd101;
vmem[4894] = 8'd116;
vmem[4895] = 8'd32;
vmem[4896] = 8'd101;
vmem[4897] = 8'd114;
vmem[4898] = 8'd111;
vmem[4899] = 8'd115;
vmem[4900] = 8'd32;
vmem[4901] = 8'd118;
vmem[4902] = 8'd101;
vmem[4903] = 8'd110;
vmem[4904] = 8'd101;
vmem[4905] = 8'd110;
vmem[4906] = 8'd97;
vmem[4907] = 8'd116;
vmem[4908] = 8'd105;
vmem[4909] = 8'd115;
vmem[4910] = 8'd32;
vmem[4911] = 8'd97;
vmem[4912] = 8'd99;
vmem[4913] = 8'd99;
vmem[4914] = 8'd117;
vmem[4915] = 8'd109;
vmem[4916] = 8'd115;
vmem[4917] = 8'd97;
vmem[4918] = 8'd110;
vmem[4919] = 8'd46;
vmem[4920] = 8'd32;
vmem[4921] = 8'd67;
vmem[4922] = 8'd117;
vmem[4923] = 8'd114;
vmem[4924] = 8'd97;
vmem[4925] = 8'd98;
vmem[4926] = 8'd105;
vmem[4927] = 8'd116;
vmem[4928] = 8'd117;
vmem[4929] = 8'd114;
vmem[4930] = 8'd32;
vmem[4931] = 8'd101;
vmem[4932] = 8'd103;
vmem[4933] = 8'd101;
vmem[4934] = 8'd116;
vmem[4935] = 8'd32;
vmem[4936] = 8'd106;
vmem[4937] = 8'd117;
vmem[4938] = 8'd115;
vmem[4939] = 8'd116;
vmem[4940] = 8'd111;
vmem[4941] = 8'd32;
vmem[4942] = 8'd110;
vmem[4943] = 8'd101;
vmem[4944] = 8'd99;
vmem[4945] = 8'd32;
vmem[4946] = 8'd108;
vmem[4947] = 8'd101;
vmem[4948] = 8'd111;
vmem[4949] = 8'd32;
vmem[4950] = 8'd118;
vmem[4951] = 8'd117;
vmem[4952] = 8'd108;
vmem[4953] = 8'd112;
vmem[4954] = 8'd117;
vmem[4955] = 8'd116;
vmem[4956] = 8'd97;
vmem[4957] = 8'd116;
vmem[4958] = 8'd101;
vmem[4959] = 8'd32;
vmem[4960] = 8'd115;
vmem[4961] = 8'd111;
vmem[4962] = 8'd108;
vmem[4963] = 8'd108;
vmem[4964] = 8'd105;
vmem[4965] = 8'd99;
vmem[4966] = 8'd105;
vmem[4967] = 8'd116;
vmem[4968] = 8'd117;
vmem[4969] = 8'd100;
vmem[4970] = 8'd105;
vmem[4971] = 8'd110;
vmem[4972] = 8'd32;
vmem[4973] = 8'd118;
vmem[4974] = 8'd101;
vmem[4975] = 8'd108;
vmem[4976] = 8'd32;
vmem[4977] = 8'd115;
vmem[4978] = 8'd101;
vmem[4979] = 8'd100;
vmem[4980] = 8'd32;
vmem[4981] = 8'd109;
vmem[4982] = 8'd105;
vmem[4983] = 8'd46;
vmem[4984] = 8'd32;
vmem[4985] = 8'd80;
vmem[4986] = 8'd104;
vmem[4987] = 8'd97;
vmem[4988] = 8'd115;
vmem[4989] = 8'd101;
vmem[4990] = 8'd108;
vmem[4991] = 8'd108;
vmem[4992] = 8'd117;
vmem[4993] = 8'd115;
vmem[4994] = 8'd32;
vmem[4995] = 8'd117;
vmem[4996] = 8'd108;
vmem[4997] = 8'd116;
vmem[4998] = 8'd114;
vmem[4999] = 8'd105;
vmem[5000] = 8'd99;
vmem[5001] = 8'd101;
vmem[5002] = 8'd115;
vmem[5003] = 8'd32;
vmem[5004] = 8'd109;
vmem[5005] = 8'd97;
vmem[5006] = 8'd103;
vmem[5007] = 8'd110;
vmem[5008] = 8'd97;
vmem[5009] = 8'd32;
vmem[5010] = 8'd99;
vmem[5011] = 8'd111;
vmem[5012] = 8'd110;
vmem[5013] = 8'd100;
vmem[5014] = 8'd105;
vmem[5015] = 8'd109;
vmem[5016] = 8'd101;
vmem[5017] = 8'd110;
vmem[5018] = 8'd116;
vmem[5019] = 8'd117;
vmem[5020] = 8'd109;
vmem[5021] = 8'd32;
vmem[5022] = 8'd108;
vmem[5023] = 8'd105;
vmem[5024] = 8'd98;
vmem[5025] = 8'd101;
vmem[5026] = 8'd114;
vmem[5027] = 8'd111;
vmem[5028] = 8'd32;
vmem[5029] = 8'd108;
vmem[5030] = 8'd97;
vmem[5031] = 8'd99;
vmem[5032] = 8'd105;
vmem[5033] = 8'd110;
vmem[5034] = 8'd105;
vmem[5035] = 8'd97;
vmem[5036] = 8'd32;
vmem[5037] = 8'd98;
vmem[5038] = 8'd105;
vmem[5039] = 8'd98;
vmem[5040] = 8'd101;
vmem[5041] = 8'd110;
vmem[5042] = 8'd100;
vmem[5043] = 8'd117;
vmem[5044] = 8'd109;
vmem[5045] = 8'd46;
vmem[5046] = 8'd32;
vmem[5047] = 8'd83;
vmem[5048] = 8'd101;
vmem[5049] = 8'd100;
vmem[5050] = 8'd32;
vmem[5051] = 8'd108;
vmem[5052] = 8'd97;
vmem[5053] = 8'd99;
vmem[5054] = 8'd117;
vmem[5055] = 8'd115;
vmem[5056] = 8'd32;
vmem[5057] = 8'd116;
vmem[5058] = 8'd117;
vmem[5059] = 8'd114;
vmem[5060] = 8'd112;
vmem[5061] = 8'd105;
vmem[5062] = 8'd115;
vmem[5063] = 8'd44;
vmem[5064] = 8'd32;
vmem[5065] = 8'd102;
vmem[5066] = 8'd101;
vmem[5067] = 8'd114;
vmem[5068] = 8'd109;
vmem[5069] = 8'd101;
vmem[5070] = 8'd110;
vmem[5071] = 8'd116;
vmem[5072] = 8'd117;
vmem[5073] = 8'd109;
vmem[5074] = 8'd32;
vmem[5075] = 8'd110;
vmem[5076] = 8'd111;
vmem[5077] = 8'd110;
vmem[5078] = 8'd32;
vmem[5079] = 8'd108;
vmem[5080] = 8'd101;
vmem[5081] = 8'd111;
vmem[5082] = 8'd32;
vmem[5083] = 8'd101;
vmem[5084] = 8'd116;
vmem[5085] = 8'd44;
vmem[5086] = 8'd32;
vmem[5087] = 8'd99;
vmem[5088] = 8'd111;
vmem[5089] = 8'd109;
vmem[5090] = 8'd109;
vmem[5091] = 8'd111;
vmem[5092] = 8'd100;
vmem[5093] = 8'd111;
vmem[5094] = 8'd32;
vmem[5095] = 8'd115;
vmem[5096] = 8'd117;
vmem[5097] = 8'd115;
vmem[5098] = 8'd99;
vmem[5099] = 8'd105;
vmem[5100] = 8'd112;
vmem[5101] = 8'd105;
vmem[5102] = 8'd116;
vmem[5103] = 8'd32;
vmem[5104] = 8'd102;
vmem[5105] = 8'd101;
vmem[5106] = 8'd108;
vmem[5107] = 8'd105;
vmem[5108] = 8'd115;
vmem[5109] = 8'd46;
vmem[5110] = 8'd32;
vmem[5111] = 8'd78;
vmem[5112] = 8'd117;
vmem[5113] = 8'd110;
vmem[5114] = 8'd99;
vmem[5115] = 8'd32;
vmem[5116] = 8'd102;
vmem[5117] = 8'd97;
vmem[5118] = 8'd117;
vmem[5119] = 8'd99;
vmem[5120] = 8'd105;
vmem[5121] = 8'd98;
vmem[5122] = 8'd117;
vmem[5123] = 8'd115;
vmem[5124] = 8'd32;
vmem[5125] = 8'd115;
vmem[5126] = 8'd101;
vmem[5127] = 8'd100;
vmem[5128] = 8'd32;
vmem[5129] = 8'd100;
vmem[5130] = 8'd117;
vmem[5131] = 8'd105;
vmem[5132] = 8'd32;
vmem[5133] = 8'd110;
vmem[5134] = 8'd101;
vmem[5135] = 8'd99;
vmem[5136] = 8'd32;
vmem[5137] = 8'd109;
vmem[5138] = 8'd111;
vmem[5139] = 8'd108;
vmem[5140] = 8'd108;
vmem[5141] = 8'd105;
vmem[5142] = 8'd115;
vmem[5143] = 8'd46;
vmem[5144] = 8'd32;
vmem[5145] = 8'd86;
vmem[5146] = 8'd105;
vmem[5147] = 8'd118;
vmem[5148] = 8'd97;
vmem[5149] = 8'd109;
vmem[5150] = 8'd117;
vmem[5151] = 8'd115;
vmem[5152] = 8'd32;
vmem[5153] = 8'd103;
vmem[5154] = 8'd114;
vmem[5155] = 8'd97;
vmem[5156] = 8'd118;
vmem[5157] = 8'd105;
vmem[5158] = 8'd100;
vmem[5159] = 8'd97;
vmem[5160] = 8'd32;
vmem[5161] = 8'd99;
vmem[5162] = 8'd111;
vmem[5163] = 8'd110;
vmem[5164] = 8'd115;
vmem[5165] = 8'd101;
vmem[5166] = 8'd113;
vmem[5167] = 8'd117;
vmem[5168] = 8'd97;
vmem[5169] = 8'd116;
vmem[5170] = 8'd32;
vmem[5171] = 8'd108;
vmem[5172] = 8'd101;
vmem[5173] = 8'd111;
vmem[5174] = 8'd46;
vmem[5175] = 8'd32;
vmem[5176] = 8'd83;
vmem[5177] = 8'd101;
vmem[5178] = 8'd100;
vmem[5179] = 8'd32;
vmem[5180] = 8'd117;
vmem[5181] = 8'd116;
vmem[5182] = 8'd32;
vmem[5183] = 8'd101;
vmem[5184] = 8'd102;
vmem[5185] = 8'd102;
vmem[5186] = 8'd105;
vmem[5187] = 8'd99;
vmem[5188] = 8'd105;
vmem[5189] = 8'd116;
vmem[5190] = 8'd117;
vmem[5191] = 8'd114;
vmem[5192] = 8'd32;
vmem[5193] = 8'd97;
vmem[5194] = 8'd114;
vmem[5195] = 8'd99;
vmem[5196] = 8'd117;
vmem[5197] = 8'd46;
vmem[5198] = 8'd32;
vmem[5199] = 8'd78;
vmem[5200] = 8'd97;
vmem[5201] = 8'd109;
vmem[5202] = 8'd32;
vmem[5203] = 8'd101;
vmem[5204] = 8'd116;
vmem[5205] = 8'd32;
vmem[5206] = 8'd101;
vmem[5207] = 8'd114;
vmem[5208] = 8'd111;
vmem[5209] = 8'd115;
vmem[5210] = 8'd32;
vmem[5211] = 8'd97;
vmem[5212] = 8'd99;
vmem[5213] = 8'd32;
vmem[5214] = 8'd101;
vmem[5215] = 8'd120;
vmem[5216] = 8'd32;
vmem[5217] = 8'd115;
vmem[5218] = 8'd111;
vmem[5219] = 8'd100;
vmem[5220] = 8'd97;
vmem[5221] = 8'd108;
vmem[5222] = 8'd101;
vmem[5223] = 8'd115;
vmem[5224] = 8'd32;
vmem[5225] = 8'd105;
vmem[5226] = 8'd110;
vmem[5227] = 8'd116;
vmem[5228] = 8'd101;
vmem[5229] = 8'd114;
vmem[5230] = 8'd100;
vmem[5231] = 8'd117;
vmem[5232] = 8'd109;
vmem[5233] = 8'd32;
vmem[5234] = 8'd101;
vmem[5235] = 8'd117;
vmem[5236] = 8'd32;
vmem[5237] = 8'd101;
vmem[5238] = 8'd103;
vmem[5239] = 8'd101;
vmem[5240] = 8'd116;
vmem[5241] = 8'd32;
vmem[5242] = 8'd108;
vmem[5243] = 8'd101;
vmem[5244] = 8'd111;
vmem[5245] = 8'd46;
vmem[5246] = 8'd32;
vmem[5247] = 8'd81;
vmem[5248] = 8'd117;
vmem[5249] = 8'd105;
vmem[5250] = 8'd115;
vmem[5251] = 8'd113;
vmem[5252] = 8'd117;
vmem[5253] = 8'd101;
vmem[5254] = 8'd32;
vmem[5255] = 8'd103;
vmem[5256] = 8'd114;
vmem[5257] = 8'd97;
vmem[5258] = 8'd118;
vmem[5259] = 8'd105;
vmem[5260] = 8'd100;
vmem[5261] = 8'd97;
vmem[5262] = 8'd32;
vmem[5263] = 8'd109;
vmem[5264] = 8'd97;
vmem[5265] = 8'd103;
vmem[5266] = 8'd110;
vmem[5267] = 8'd97;
vmem[5268] = 8'd32;
vmem[5269] = 8'd108;
vmem[5270] = 8'd101;
vmem[5271] = 8'd111;
vmem[5272] = 8'd44;
vmem[5273] = 8'd32;
vmem[5274] = 8'd101;
vmem[5275] = 8'd116;
vmem[5276] = 8'd32;
vmem[5277] = 8'd118;
vmem[5278] = 8'd117;
vmem[5279] = 8'd108;
vmem[5280] = 8'd112;
vmem[5281] = 8'd117;
vmem[5282] = 8'd116;
vmem[5283] = 8'd97;
vmem[5284] = 8'd116;
vmem[5285] = 8'd101;
vmem[5286] = 8'd32;
vmem[5287] = 8'd110;
vmem[5288] = 8'd105;
vmem[5289] = 8'd115;
vmem[5290] = 8'd105;
vmem[5291] = 8'd32;
vmem[5292] = 8'd98;
vmem[5293] = 8'd108;
vmem[5294] = 8'd97;
vmem[5295] = 8'd110;
vmem[5296] = 8'd100;
vmem[5297] = 8'd105;
vmem[5298] = 8'd116;
vmem[5299] = 8'd32;
vmem[5300] = 8'd113;
vmem[5301] = 8'd117;
vmem[5302] = 8'd105;
vmem[5303] = 8'd115;
vmem[5304] = 8'd46;
vmem[5305] = 8'd32;
vmem[5306] = 8'd68;
vmem[5307] = 8'd117;
vmem[5308] = 8'd105;
vmem[5309] = 8'd115;
vmem[5310] = 8'd32;
vmem[5311] = 8'd101;
vmem[5312] = 8'd103;
vmem[5313] = 8'd101;
vmem[5314] = 8'd116;
vmem[5315] = 8'd32;
vmem[5316] = 8'd112;
vmem[5317] = 8'd111;
vmem[5318] = 8'd114;
vmem[5319] = 8'd116;
vmem[5320] = 8'd116;
vmem[5321] = 8'd105;
vmem[5322] = 8'd116;
vmem[5323] = 8'd111;
vmem[5324] = 8'd114;
vmem[5325] = 8'd32;
vmem[5326] = 8'd110;
vmem[5327] = 8'd117;
vmem[5328] = 8'd108;
vmem[5329] = 8'd108;
vmem[5330] = 8'd97;
vmem[5331] = 8'd46;
vmem[5332] = 8'd32;
vmem[5333] = 8'd67;
vmem[5334] = 8'd114;
vmem[5335] = 8'd97;
vmem[5336] = 8'd115;
vmem[5337] = 8'd32;
vmem[5338] = 8'd109;
vmem[5339] = 8'd97;
vmem[5340] = 8'd108;
vmem[5341] = 8'd101;
vmem[5342] = 8'd115;
vmem[5343] = 8'd117;
vmem[5344] = 8'd97;
vmem[5345] = 8'd100;
vmem[5346] = 8'd97;
vmem[5347] = 8'd32;
vmem[5348] = 8'd112;
vmem[5349] = 8'd108;
vmem[5350] = 8'd97;
vmem[5351] = 8'd99;
vmem[5352] = 8'd101;
vmem[5353] = 8'd114;
vmem[5354] = 8'd97;
vmem[5355] = 8'd116;
vmem[5356] = 8'd32;
vmem[5357] = 8'd110;
vmem[5358] = 8'd117;
vmem[5359] = 8'd110;
vmem[5360] = 8'd99;
vmem[5361] = 8'd32;
vmem[5362] = 8'd101;
vmem[5363] = 8'd103;
vmem[5364] = 8'd101;
vmem[5365] = 8'd116;
vmem[5366] = 8'd32;
vmem[5367] = 8'd100;
vmem[5368] = 8'd97;
vmem[5369] = 8'd112;
vmem[5370] = 8'd105;
vmem[5371] = 8'd98;
vmem[5372] = 8'd117;
vmem[5373] = 8'd115;
vmem[5374] = 8'd46;
vmem[5375] = 8'd32;
vmem[5376] = 8'd65;
vmem[5377] = 8'd108;
vmem[5378] = 8'd105;
vmem[5379] = 8'd113;
vmem[5380] = 8'd117;
vmem[5381] = 8'd97;
vmem[5382] = 8'd109;
vmem[5383] = 8'd32;
vmem[5384] = 8'd117;
vmem[5385] = 8'd108;
vmem[5386] = 8'd116;
vmem[5387] = 8'd114;
vmem[5388] = 8'd105;
vmem[5389] = 8'd99;
vmem[5390] = 8'd101;
vmem[5391] = 8'd115;
vmem[5392] = 8'd32;
vmem[5393] = 8'd112;
vmem[5394] = 8'd117;
vmem[5395] = 8'd108;
vmem[5396] = 8'd118;
vmem[5397] = 8'd105;
vmem[5398] = 8'd110;
vmem[5399] = 8'd97;
vmem[5400] = 8'd114;
vmem[5401] = 8'd32;
vmem[5402] = 8'd118;
vmem[5403] = 8'd97;
vmem[5404] = 8'd114;
vmem[5405] = 8'd105;
vmem[5406] = 8'd117;
vmem[5407] = 8'd115;
vmem[5408] = 8'd46;
vmem[5409] = 8'd32;
vmem[5410] = 8'd80;
vmem[5411] = 8'd114;
vmem[5412] = 8'd111;
vmem[5413] = 8'd105;
vmem[5414] = 8'd110;
vmem[5415] = 8'd32;
vmem[5416] = 8'd108;
vmem[5417] = 8'd97;
vmem[5418] = 8'd111;
vmem[5419] = 8'd114;
vmem[5420] = 8'd101;
vmem[5421] = 8'd101;
vmem[5422] = 8'd116;
vmem[5423] = 8'd32;
vmem[5424] = 8'd108;
vmem[5425] = 8'd101;
vmem[5426] = 8'd99;
vmem[5427] = 8'd116;
vmem[5428] = 8'd117;
vmem[5429] = 8'd115;
vmem[5430] = 8'd32;
vmem[5431] = 8'd101;
vmem[5432] = 8'd117;
vmem[5433] = 8'd32;
vmem[5434] = 8'd102;
vmem[5435] = 8'd105;
vmem[5436] = 8'd110;
vmem[5437] = 8'd105;
vmem[5438] = 8'd98;
vmem[5439] = 8'd117;
vmem[5440] = 8'd115;
vmem[5441] = 8'd32;
vmem[5442] = 8'd99;
vmem[5443] = 8'd111;
vmem[5444] = 8'd110;
vmem[5445] = 8'd115;
vmem[5446] = 8'd101;
vmem[5447] = 8'd99;
vmem[5448] = 8'd116;
vmem[5449] = 8'd101;
vmem[5450] = 8'd116;
vmem[5451] = 8'd117;
vmem[5452] = 8'd114;
vmem[5453] = 8'd46;
vmem[5454] = 8'd32;
vmem[5455] = 8'd65;
vmem[5456] = 8'd108;
vmem[5457] = 8'd105;
vmem[5458] = 8'd113;
vmem[5459] = 8'd117;
vmem[5460] = 8'd97;
vmem[5461] = 8'd109;
vmem[5462] = 8'd32;
vmem[5463] = 8'd101;
vmem[5464] = 8'd114;
vmem[5465] = 8'd97;
vmem[5466] = 8'd116;
vmem[5467] = 8'd32;
vmem[5468] = 8'd118;
vmem[5469] = 8'd111;
vmem[5470] = 8'd108;
vmem[5471] = 8'd117;
vmem[5472] = 8'd116;
vmem[5473] = 8'd112;
vmem[5474] = 8'd97;
vmem[5475] = 8'd116;
vmem[5476] = 8'd46;
vmem[5477] = 8'd32;
vmem[5478] = 8'd73;
vmem[5479] = 8'd110;
vmem[5480] = 8'd32;
vmem[5481] = 8'd99;
vmem[5482] = 8'd117;
vmem[5483] = 8'd114;
vmem[5484] = 8'd115;
vmem[5485] = 8'd117;
vmem[5486] = 8'd115;
vmem[5487] = 8'd32;
vmem[5488] = 8'd117;
vmem[5489] = 8'd114;
vmem[5490] = 8'd110;
vmem[5491] = 8'd97;
vmem[5492] = 8'd32;
vmem[5493] = 8'd101;
vmem[5494] = 8'd117;
vmem[5495] = 8'd32;
vmem[5496] = 8'd109;
vmem[5497] = 8'd97;
vmem[5498] = 8'd103;
vmem[5499] = 8'd110;
vmem[5500] = 8'd97;
vmem[5501] = 8'd32;
vmem[5502] = 8'd108;
vmem[5503] = 8'd97;
vmem[5504] = 8'd99;
vmem[5505] = 8'd105;
vmem[5506] = 8'd110;
vmem[5507] = 8'd105;
vmem[5508] = 8'd97;
vmem[5509] = 8'd44;
vmem[5510] = 8'd32;
vmem[5511] = 8'd97;
vmem[5512] = 8'd99;
vmem[5513] = 8'd32;
vmem[5514] = 8'd117;
vmem[5515] = 8'd108;
vmem[5516] = 8'd108;
vmem[5517] = 8'd97;
vmem[5518] = 8'd109;
vmem[5519] = 8'd99;
vmem[5520] = 8'd111;
vmem[5521] = 8'd114;
vmem[5522] = 8'd112;
vmem[5523] = 8'd101;
vmem[5524] = 8'd114;
vmem[5525] = 8'd32;
vmem[5526] = 8'd108;
vmem[5527] = 8'd105;
vmem[5528] = 8'd103;
vmem[5529] = 8'd117;
vmem[5530] = 8'd108;
vmem[5531] = 8'd97;
vmem[5532] = 8'd32;
vmem[5533] = 8'd98;
vmem[5534] = 8'd108;
vmem[5535] = 8'd97;
vmem[5536] = 8'd110;
vmem[5537] = 8'd100;
vmem[5538] = 8'd105;
vmem[5539] = 8'd116;
vmem[5540] = 8'd46;
vmem[5541] = 8'd32;
vmem[5542] = 8'd85;
vmem[5543] = 8'd116;
vmem[5544] = 8'd32;
vmem[5545] = 8'd112;
vmem[5546] = 8'd101;
vmem[5547] = 8'd108;
vmem[5548] = 8'd108;
vmem[5549] = 8'd101;
vmem[5550] = 8'd110;
vmem[5551] = 8'd116;
vmem[5552] = 8'd101;
vmem[5553] = 8'd115;
vmem[5554] = 8'd113;
vmem[5555] = 8'd117;
vmem[5556] = 8'd101;
vmem[5557] = 8'd32;
vmem[5558] = 8'd97;
vmem[5559] = 8'd117;
vmem[5560] = 8'd103;
vmem[5561] = 8'd117;
vmem[5562] = 8'd101;
vmem[5563] = 8'd32;
vmem[5564] = 8'd101;
vmem[5565] = 8'd110;
vmem[5566] = 8'd105;
vmem[5567] = 8'd109;
vmem[5568] = 8'd44;
vmem[5569] = 8'd32;
vmem[5570] = 8'd101;
vmem[5571] = 8'd103;
vmem[5572] = 8'd101;
vmem[5573] = 8'd116;
vmem[5574] = 8'd32;
vmem[5575] = 8'd102;
vmem[5576] = 8'd97;
vmem[5577] = 8'd117;
vmem[5578] = 8'd99;
vmem[5579] = 8'd105;
vmem[5580] = 8'd98;
vmem[5581] = 8'd117;
vmem[5582] = 8'd115;
vmem[5583] = 8'd32;
vmem[5584] = 8'd110;
vmem[5585] = 8'd101;
vmem[5586] = 8'd113;
vmem[5587] = 8'd117;
vmem[5588] = 8'd101;
vmem[5589] = 8'd32;
vmem[5590] = 8'd102;
vmem[5591] = 8'd101;
vmem[5592] = 8'd114;
vmem[5593] = 8'd109;
vmem[5594] = 8'd101;
vmem[5595] = 8'd110;
vmem[5596] = 8'd116;
vmem[5597] = 8'd117;
vmem[5598] = 8'd109;
vmem[5599] = 8'd32;
vmem[5600] = 8'd97;
vmem[5601] = 8'd99;
vmem[5602] = 8'd46;
vmem[5603] = 8'd32;
vmem[5604] = 8'd83;
vmem[5605] = 8'd117;
vmem[5606] = 8'd115;
vmem[5607] = 8'd112;
vmem[5608] = 8'd101;
vmem[5609] = 8'd110;
vmem[5610] = 8'd100;
vmem[5611] = 8'd105;
vmem[5612] = 8'd115;
vmem[5613] = 8'd115;
vmem[5614] = 8'd101;
vmem[5615] = 8'd32;
vmem[5616] = 8'd97;
vmem[5617] = 8'd99;
vmem[5618] = 8'd32;
vmem[5619] = 8'd99;
vmem[5620] = 8'd111;
vmem[5621] = 8'd110;
vmem[5622] = 8'd115;
vmem[5623] = 8'd101;
vmem[5624] = 8'd99;
vmem[5625] = 8'd116;
vmem[5626] = 8'd101;
vmem[5627] = 8'd116;
vmem[5628] = 8'd117;
vmem[5629] = 8'd114;
vmem[5630] = 8'd32;
vmem[5631] = 8'd117;
vmem[5632] = 8'd114;
vmem[5633] = 8'd110;
vmem[5634] = 8'd97;
vmem[5635] = 8'd46;
vmem[5636] = 8'd32;
vmem[5637] = 8'd80;
vmem[5638] = 8'd114;
vmem[5639] = 8'd97;
vmem[5640] = 8'd101;
vmem[5641] = 8'd115;
vmem[5642] = 8'd101;
vmem[5643] = 8'd110;
vmem[5644] = 8'd116;
vmem[5645] = 8'd32;
vmem[5646] = 8'd115;
vmem[5647] = 8'd101;
vmem[5648] = 8'd109;
vmem[5649] = 8'd112;
vmem[5650] = 8'd101;
vmem[5651] = 8'd114;
vmem[5652] = 8'd32;
vmem[5653] = 8'd118;
vmem[5654] = 8'd101;
vmem[5655] = 8'd108;
vmem[5656] = 8'd105;
vmem[5657] = 8'd116;
vmem[5658] = 8'd32;
vmem[5659] = 8'd105;
vmem[5660] = 8'd110;
vmem[5661] = 8'd32;
vmem[5662] = 8'd100;
vmem[5663] = 8'd105;
vmem[5664] = 8'd97;
vmem[5665] = 8'd109;
vmem[5666] = 8'd32;
vmem[5667] = 8'd99;
vmem[5668] = 8'd117;
vmem[5669] = 8'd114;
vmem[5670] = 8'd115;
vmem[5671] = 8'd117;
vmem[5672] = 8'd115;
vmem[5673] = 8'd32;
vmem[5674] = 8'd112;
vmem[5675] = 8'd104;
vmem[5676] = 8'd97;
vmem[5677] = 8'd114;
vmem[5678] = 8'd101;
vmem[5679] = 8'd116;
vmem[5680] = 8'd114;
vmem[5681] = 8'd97;
vmem[5682] = 8'd46;
vmem[5683] = 8'd32;
vmem[5684] = 8'd65;
vmem[5685] = 8'd108;
vmem[5686] = 8'd105;
vmem[5687] = 8'd113;
vmem[5688] = 8'd117;
vmem[5689] = 8'd97;
vmem[5690] = 8'd109;
vmem[5691] = 8'd32;
vmem[5692] = 8'd101;
vmem[5693] = 8'd114;
vmem[5694] = 8'd97;
vmem[5695] = 8'd116;
vmem[5696] = 8'd32;
vmem[5697] = 8'd118;
vmem[5698] = 8'd111;
vmem[5699] = 8'd108;
vmem[5700] = 8'd117;
vmem[5701] = 8'd116;
vmem[5702] = 8'd112;
vmem[5703] = 8'd97;
vmem[5704] = 8'd116;
vmem[5705] = 8'd46;
vmem[5706] = 8'd32;
vmem[5707] = 8'd77;
vmem[5708] = 8'd111;
vmem[5709] = 8'd114;
vmem[5710] = 8'd98;
vmem[5711] = 8'd105;
vmem[5712] = 8'd32;
vmem[5713] = 8'd115;
vmem[5714] = 8'd105;
vmem[5715] = 8'd116;
vmem[5716] = 8'd32;
vmem[5717] = 8'd97;
vmem[5718] = 8'd109;
vmem[5719] = 8'd101;
vmem[5720] = 8'd116;
vmem[5721] = 8'd32;
vmem[5722] = 8'd115;
vmem[5723] = 8'd111;
vmem[5724] = 8'd108;
vmem[5725] = 8'd108;
vmem[5726] = 8'd105;
vmem[5727] = 8'd99;
vmem[5728] = 8'd105;
vmem[5729] = 8'd116;
vmem[5730] = 8'd117;
vmem[5731] = 8'd100;
vmem[5732] = 8'd105;
vmem[5733] = 8'd110;
vmem[5734] = 8'd32;
vmem[5735] = 8'd111;
vmem[5736] = 8'd114;
vmem[5737] = 8'd99;
vmem[5738] = 8'd105;
vmem[5739] = 8'd44;
vmem[5740] = 8'd32;
vmem[5741] = 8'd101;
vmem[5742] = 8'd103;
vmem[5743] = 8'd101;
vmem[5744] = 8'd116;
vmem[5745] = 8'd32;
vmem[5746] = 8'd99;
vmem[5747] = 8'd111;
vmem[5748] = 8'd110;
vmem[5749] = 8'd115;
vmem[5750] = 8'd101;
vmem[5751] = 8'd99;
vmem[5752] = 8'd116;
vmem[5753] = 8'd101;
vmem[5754] = 8'd116;
vmem[5755] = 8'd117;
vmem[5756] = 8'd114;
vmem[5757] = 8'd32;
vmem[5758] = 8'd102;
vmem[5759] = 8'd101;
vmem[5760] = 8'd108;
vmem[5761] = 8'd105;
vmem[5762] = 8'd115;
vmem[5763] = 8'd46;
vmem[5764] = 8'd32;
vmem[5765] = 8'd78;
vmem[5766] = 8'd97;
vmem[5767] = 8'd109;
vmem[5768] = 8'd32;
vmem[5769] = 8'd105;
vmem[5770] = 8'd100;
vmem[5771] = 8'd32;
vmem[5772] = 8'd108;
vmem[5773] = 8'd101;
vmem[5774] = 8'd99;
vmem[5775] = 8'd116;
vmem[5776] = 8'd117;
vmem[5777] = 8'd115;
vmem[5778] = 8'd32;
vmem[5779] = 8'd118;
vmem[5780] = 8'd101;
vmem[5781] = 8'd108;
vmem[5782] = 8'd32;
vmem[5783] = 8'd108;
vmem[5784] = 8'd101;
vmem[5785] = 8'd111;
vmem[5786] = 8'd32;
vmem[5787] = 8'd108;
vmem[5788] = 8'd117;
vmem[5789] = 8'd99;
vmem[5790] = 8'd116;
vmem[5791] = 8'd117;
vmem[5792] = 8'd115;
vmem[5793] = 8'd32;
vmem[5794] = 8'd109;
vmem[5795] = 8'd111;
vmem[5796] = 8'd108;
vmem[5797] = 8'd108;
vmem[5798] = 8'd105;
vmem[5799] = 8'd115;
vmem[5800] = 8'd32;
vmem[5801] = 8'd101;
vmem[5802] = 8'd116;
vmem[5803] = 8'd32;
vmem[5804] = 8'd118;
vmem[5805] = 8'd101;
vmem[5806] = 8'd108;
vmem[5807] = 8'd32;
vmem[5808] = 8'd100;
vmem[5809] = 8'd117;
vmem[5810] = 8'd105;
vmem[5811] = 8'd46;
vmem[5812] = 8'd32;
vmem[5813] = 8'd78;
vmem[5814] = 8'd117;
vmem[5815] = 8'd108;
vmem[5816] = 8'd108;
vmem[5817] = 8'd97;
vmem[5818] = 8'd109;
vmem[5819] = 8'd32;
vmem[5820] = 8'd101;
vmem[5821] = 8'd120;
vmem[5822] = 8'd32;
vmem[5823] = 8'd112;
vmem[5824] = 8'd117;
vmem[5825] = 8'd114;
vmem[5826] = 8'd117;
vmem[5827] = 8'd115;
vmem[5828] = 8'd44;
vmem[5829] = 8'd32;
vmem[5830] = 8'd116;
vmem[5831] = 8'd105;
vmem[5832] = 8'd110;
vmem[5833] = 8'd99;
vmem[5834] = 8'd105;
vmem[5835] = 8'd100;
vmem[5836] = 8'd117;
vmem[5837] = 8'd110;
vmem[5838] = 8'd116;
vmem[5839] = 8'd32;
vmem[5840] = 8'd118;
vmem[5841] = 8'd101;
vmem[5842] = 8'd108;
vmem[5843] = 8'd32;
vmem[5844] = 8'd109;
vmem[5845] = 8'd105;
vmem[5846] = 8'd32;
vmem[5847] = 8'd110;
vmem[5848] = 8'd111;
vmem[5849] = 8'd110;
vmem[5850] = 8'd44;
vmem[5851] = 8'd32;
vmem[5852] = 8'd112;
vmem[5853] = 8'd114;
vmem[5854] = 8'd101;
vmem[5855] = 8'd116;
vmem[5856] = 8'd105;
vmem[5857] = 8'd117;
vmem[5858] = 8'd109;
vmem[5859] = 8'd32;
vmem[5860] = 8'd118;
vmem[5861] = 8'd101;
vmem[5862] = 8'd110;
vmem[5863] = 8'd101;
vmem[5864] = 8'd110;
vmem[5865] = 8'd97;
vmem[5866] = 8'd116;
vmem[5867] = 8'd105;
vmem[5868] = 8'd115;
vmem[5869] = 8'd32;
vmem[5870] = 8'd105;
vmem[5871] = 8'd112;
vmem[5872] = 8'd115;
vmem[5873] = 8'd117;
vmem[5874] = 8'd109;
vmem[5875] = 8'd46;
vmem[5876] = 8'd32;
vmem[5877] = 8'd77;
vmem[5878] = 8'd97;
vmem[5879] = 8'd101;
vmem[5880] = 8'd99;
vmem[5881] = 8'd101;
vmem[5882] = 8'd110;
vmem[5883] = 8'd97;
vmem[5884] = 8'd115;
vmem[5885] = 8'd32;
vmem[5886] = 8'd101;
vmem[5887] = 8'd103;
vmem[5888] = 8'd101;
vmem[5889] = 8'd116;
vmem[5890] = 8'd32;
vmem[5891] = 8'd109;
vmem[5892] = 8'd97;
vmem[5893] = 8'd108;
vmem[5894] = 8'd101;
vmem[5895] = 8'd115;
vmem[5896] = 8'd117;
vmem[5897] = 8'd97;
vmem[5898] = 8'd100;
vmem[5899] = 8'd97;
vmem[5900] = 8'd32;
vmem[5901] = 8'd115;
vmem[5902] = 8'd101;
vmem[5903] = 8'd109;
vmem[5904] = 8'd46;
vmem[5905] = 8'd32;
vmem[5906] = 8'd80;
vmem[5907] = 8'd114;
vmem[5908] = 8'd97;
vmem[5909] = 8'd101;
vmem[5910] = 8'd115;
vmem[5911] = 8'd101;
vmem[5912] = 8'd110;
vmem[5913] = 8'd116;
vmem[5914] = 8'd32;
vmem[5915] = 8'd101;
vmem[5916] = 8'd108;
vmem[5917] = 8'd101;
vmem[5918] = 8'd109;
vmem[5919] = 8'd101;
vmem[5920] = 8'd110;
vmem[5921] = 8'd116;
vmem[5922] = 8'd117;
vmem[5923] = 8'd109;
vmem[5924] = 8'd32;
vmem[5925] = 8'd115;
vmem[5926] = 8'd99;
vmem[5927] = 8'd101;
vmem[5928] = 8'd108;
vmem[5929] = 8'd101;
vmem[5930] = 8'd114;
vmem[5931] = 8'd105;
vmem[5932] = 8'd115;
vmem[5933] = 8'd113;
vmem[5934] = 8'd117;
vmem[5935] = 8'd101;
vmem[5936] = 8'd32;
vmem[5937] = 8'd118;
vmem[5938] = 8'd101;
vmem[5939] = 8'd108;
vmem[5940] = 8'd105;
vmem[5941] = 8'd116;
vmem[5942] = 8'd44;
vmem[5943] = 8'd32;
vmem[5944] = 8'd105;
vmem[5945] = 8'd110;
vmem[5946] = 8'd32;
vmem[5947] = 8'd101;
vmem[5948] = 8'd117;
vmem[5949] = 8'd105;
vmem[5950] = 8'd115;
vmem[5951] = 8'd109;
vmem[5952] = 8'd111;
vmem[5953] = 8'd100;
vmem[5954] = 8'd32;
vmem[5955] = 8'd118;
vmem[5956] = 8'd101;
vmem[5957] = 8'd108;
vmem[5958] = 8'd105;
vmem[5959] = 8'd116;
vmem[5960] = 8'd32;
vmem[5961] = 8'd116;
vmem[5962] = 8'd114;
vmem[5963] = 8'd105;
vmem[5964] = 8'd115;
vmem[5965] = 8'd116;
vmem[5966] = 8'd105;
vmem[5967] = 8'd113;
vmem[5968] = 8'd117;
vmem[5969] = 8'd101;
vmem[5970] = 8'd32;
vmem[5971] = 8'd105;
vmem[5972] = 8'd109;
vmem[5973] = 8'd112;
vmem[5974] = 8'd101;
vmem[5975] = 8'd114;
vmem[5976] = 8'd100;
vmem[5977] = 8'd105;
vmem[5978] = 8'd101;
vmem[5979] = 8'd116;
vmem[5980] = 8'd46;
vmem[5981] = 8'd32;
vmem[5982] = 8'd78;
vmem[5983] = 8'd97;
vmem[5984] = 8'd109;
vmem[5985] = 8'd32;
vmem[5986] = 8'd116;
vmem[5987] = 8'd101;
vmem[5988] = 8'd109;
vmem[5989] = 8'd112;
vmem[5990] = 8'd111;
vmem[5991] = 8'd114;
vmem[5992] = 8'd44;
vmem[5993] = 8'd32;
vmem[5994] = 8'd108;
vmem[5995] = 8'd105;
vmem[5996] = 8'd98;
vmem[5997] = 8'd101;
vmem[5998] = 8'd114;
vmem[5999] = 8'd111;
vmem[6000] = 8'd32;
vmem[6001] = 8'd103;
vmem[6002] = 8'd114;
vmem[6003] = 8'd97;
vmem[6004] = 8'd118;
vmem[6005] = 8'd105;
vmem[6006] = 8'd100;
vmem[6007] = 8'd97;
vmem[6008] = 8'd32;
vmem[6009] = 8'd116;
vmem[6010] = 8'd114;
vmem[6011] = 8'd105;
vmem[6012] = 8'd115;
vmem[6013] = 8'd116;
vmem[6014] = 8'd105;
vmem[6015] = 8'd113;
vmem[6016] = 8'd117;
vmem[6017] = 8'd101;
vmem[6018] = 8'd32;
vmem[6019] = 8'd111;
vmem[6020] = 8'd114;
vmem[6021] = 8'd110;
vmem[6022] = 8'd97;
vmem[6023] = 8'd114;
vmem[6024] = 8'd101;
vmem[6025] = 8'd44;
vmem[6026] = 8'd32;
vmem[6027] = 8'd117;
vmem[6028] = 8'd114;
vmem[6029] = 8'd110;
vmem[6030] = 8'd97;
vmem[6031] = 8'd32;
vmem[6032] = 8'd109;
vmem[6033] = 8'd97;
vmem[6034] = 8'd103;
vmem[6035] = 8'd110;
vmem[6036] = 8'd97;
vmem[6037] = 8'd32;
vmem[6038] = 8'd118;
vmem[6039] = 8'd105;
vmem[6040] = 8'd118;
vmem[6041] = 8'd101;
vmem[6042] = 8'd114;
vmem[6043] = 8'd114;
vmem[6044] = 8'd97;
vmem[6045] = 8'd32;
vmem[6046] = 8'd100;
vmem[6047] = 8'd117;
vmem[6048] = 8'd105;
vmem[6049] = 8'd44;
vmem[6050] = 8'd32;
vmem[6051] = 8'd105;
vmem[6052] = 8'd110;
vmem[6053] = 8'd116;
vmem[6054] = 8'd101;
vmem[6055] = 8'd114;
vmem[6056] = 8'd100;
vmem[6057] = 8'd117;
vmem[6058] = 8'd109;
vmem[6059] = 8'd32;
vmem[6060] = 8'd99;
vmem[6061] = 8'd111;
vmem[6062] = 8'd110;
vmem[6063] = 8'd103;
vmem[6064] = 8'd117;
vmem[6065] = 8'd101;
vmem[6066] = 8'd32;
vmem[6067] = 8'd112;
vmem[6068] = 8'd117;
vmem[6069] = 8'd114;
vmem[6070] = 8'd117;
vmem[6071] = 8'd115;
vmem[6072] = 8'd32;
vmem[6073] = 8'd116;
vmem[6074] = 8'd111;
vmem[6075] = 8'd114;
vmem[6076] = 8'd116;
vmem[6077] = 8'd111;
vmem[6078] = 8'd114;
vmem[6079] = 8'd32;
vmem[6080] = 8'd102;
vmem[6081] = 8'd105;
vmem[6082] = 8'd110;
vmem[6083] = 8'd105;
vmem[6084] = 8'd98;
vmem[6085] = 8'd117;
vmem[6086] = 8'd115;
vmem[6087] = 8'd32;
vmem[6088] = 8'd108;
vmem[6089] = 8'd101;
vmem[6090] = 8'd99;
vmem[6091] = 8'd116;
vmem[6092] = 8'd117;
vmem[6093] = 8'd115;
vmem[6094] = 8'd46;
vmem[6095] = 8'd32;
vmem[6096] = 8'd77;
vmem[6097] = 8'd97;
vmem[6098] = 8'd101;
vmem[6099] = 8'd99;
vmem[6100] = 8'd101;
vmem[6101] = 8'd110;
vmem[6102] = 8'd97;
vmem[6103] = 8'd115;
vmem[6104] = 8'd32;
vmem[6105] = 8'd109;
vmem[6106] = 8'd97;
vmem[6107] = 8'd108;
vmem[6108] = 8'd101;
vmem[6109] = 8'd115;
vmem[6110] = 8'd117;
vmem[6111] = 8'd97;
vmem[6112] = 8'd100;
vmem[6113] = 8'd97;
vmem[6114] = 8'd32;
vmem[6115] = 8'd97;
vmem[6116] = 8'd99;
vmem[6117] = 8'd32;
vmem[6118] = 8'd110;
vmem[6119] = 8'd105;
vmem[6120] = 8'd98;
vmem[6121] = 8'd104;
vmem[6122] = 8'd32;
vmem[6123] = 8'd115;
vmem[6124] = 8'd105;
vmem[6125] = 8'd116;
vmem[6126] = 8'd32;
vmem[6127] = 8'd97;
vmem[6128] = 8'd109;
vmem[6129] = 8'd101;
vmem[6130] = 8'd116;
vmem[6131] = 8'd32;
vmem[6132] = 8'd118;
vmem[6133] = 8'd117;
vmem[6134] = 8'd108;
vmem[6135] = 8'd112;
vmem[6136] = 8'd117;
vmem[6137] = 8'd116;
vmem[6138] = 8'd97;
vmem[6139] = 8'd116;
vmem[6140] = 8'd101;
vmem[6141] = 8'd46;
vmem[6142] = 8'd32;
vmem[6143] = 8'd86;
vmem[6144] = 8'd101;
vmem[6145] = 8'd115;
vmem[6146] = 8'd116;
vmem[6147] = 8'd105;
vmem[6148] = 8'd98;
vmem[6149] = 8'd117;
vmem[6150] = 8'd108;
vmem[6151] = 8'd117;
vmem[6152] = 8'd109;
vmem[6153] = 8'd32;
vmem[6154] = 8'd118;
vmem[6155] = 8'd105;
vmem[6156] = 8'd116;
vmem[6157] = 8'd97;
vmem[6158] = 8'd101;
vmem[6159] = 8'd32;
vmem[6160] = 8'd110;
vmem[6161] = 8'd105;
vmem[6162] = 8'd115;
vmem[6163] = 8'd105;
vmem[6164] = 8'd32;
vmem[6165] = 8'd110;
vmem[6166] = 8'd105;
vmem[6167] = 8'd115;
vmem[6168] = 8'd105;
vmem[6169] = 8'd46;
vmem[6170] = 8'd32;
vmem[6171] = 8'd67;
vmem[6172] = 8'd114;
vmem[6173] = 8'd97;
vmem[6174] = 8'd115;
vmem[6175] = 8'd32;
vmem[6176] = 8'd117;
vmem[6177] = 8'd108;
vmem[6178] = 8'd116;
vmem[6179] = 8'd114;
vmem[6180] = 8'd105;
vmem[6181] = 8'd99;
vmem[6182] = 8'd101;
vmem[6183] = 8'd115;
vmem[6184] = 8'd32;
vmem[6185] = 8'd113;
vmem[6186] = 8'd117;
vmem[6187] = 8'd105;
vmem[6188] = 8'd115;
vmem[6189] = 8'd32;
vmem[6190] = 8'd100;
vmem[6191] = 8'd111;
vmem[6192] = 8'd108;
vmem[6193] = 8'd111;
vmem[6194] = 8'd114;
vmem[6195] = 8'd32;
vmem[6196] = 8'd110;
vmem[6197] = 8'd111;
vmem[6198] = 8'd110;
vmem[6199] = 8'd32;
vmem[6200] = 8'd97;
vmem[6201] = 8'd108;
vmem[6202] = 8'd105;
vmem[6203] = 8'd113;
vmem[6204] = 8'd117;
vmem[6205] = 8'd101;
vmem[6206] = 8'd116;
vmem[6207] = 8'd46;
vmem[6208] = 8'd32;
vmem[6209] = 8'd68;
vmem[6210] = 8'd117;
vmem[6211] = 8'd105;
vmem[6212] = 8'd115;
vmem[6213] = 8'd32;
vmem[6214] = 8'd100;
vmem[6215] = 8'd105;
vmem[6216] = 8'd97;
vmem[6217] = 8'd109;
vmem[6218] = 8'd32;
vmem[6219] = 8'd113;
vmem[6220] = 8'd117;
vmem[6221] = 8'd97;
vmem[6222] = 8'd109;
vmem[6223] = 8'd44;
vmem[6224] = 8'd32;
vmem[6225] = 8'd102;
vmem[6226] = 8'd105;
vmem[6227] = 8'd110;
vmem[6228] = 8'd105;
vmem[6229] = 8'd98;
vmem[6230] = 8'd117;
vmem[6231] = 8'd115;
vmem[6232] = 8'd32;
vmem[6233] = 8'd105;
vmem[6234] = 8'd110;
vmem[6235] = 8'd32;
vmem[6236] = 8'd102;
vmem[6237] = 8'd101;
vmem[6238] = 8'd108;
vmem[6239] = 8'd105;
vmem[6240] = 8'd115;
vmem[6241] = 8'd32;
vmem[6242] = 8'd110;
vmem[6243] = 8'd101;
vmem[6244] = 8'd99;
vmem[6245] = 8'd44;
vmem[6246] = 8'd32;
vmem[6247] = 8'd117;
vmem[6248] = 8'd108;
vmem[6249] = 8'd116;
vmem[6250] = 8'd114;
vmem[6251] = 8'd105;
vmem[6252] = 8'd99;
vmem[6253] = 8'd105;
vmem[6254] = 8'd101;
vmem[6255] = 8'd115;
vmem[6256] = 8'd32;
vmem[6257] = 8'd109;
vmem[6258] = 8'd111;
vmem[6259] = 8'd108;
vmem[6260] = 8'd101;
vmem[6261] = 8'd115;
vmem[6262] = 8'd116;
vmem[6263] = 8'd105;
vmem[6264] = 8'd101;
vmem[6265] = 8'd32;
vmem[6266] = 8'd108;
vmem[6267] = 8'd105;
vmem[6268] = 8'd103;
vmem[6269] = 8'd117;
vmem[6270] = 8'd108;
vmem[6271] = 8'd97;
vmem[6272] = 8'd46;
vmem[6273] = 8'd32;
vmem[6274] = 8'd67;
vmem[6275] = 8'd117;
vmem[6276] = 8'd114;
vmem[6277] = 8'd97;
vmem[6278] = 8'd98;
vmem[6279] = 8'd105;
vmem[6280] = 8'd116;
vmem[6281] = 8'd117;
vmem[6282] = 8'd114;
vmem[6283] = 8'd32;
vmem[6284] = 8'd110;
vmem[6285] = 8'd105;
vmem[6286] = 8'd115;
vmem[6287] = 8'd105;
vmem[6288] = 8'd32;
vmem[6289] = 8'd97;
vmem[6290] = 8'd114;
vmem[6291] = 8'd99;
vmem[6292] = 8'd117;
vmem[6293] = 8'd44;
vmem[6294] = 8'd32;
vmem[6295] = 8'd97;
vmem[6296] = 8'd99;
vmem[6297] = 8'd99;
vmem[6298] = 8'd117;
vmem[6299] = 8'd109;
vmem[6300] = 8'd115;
vmem[6301] = 8'd97;
vmem[6302] = 8'd110;
vmem[6303] = 8'd32;
vmem[6304] = 8'd113;
vmem[6305] = 8'd117;
vmem[6306] = 8'd105;
vmem[6307] = 8'd115;
vmem[6308] = 8'd32;
vmem[6309] = 8'd99;
vmem[6310] = 8'd111;
vmem[6311] = 8'd110;
vmem[6312] = 8'd100;
vmem[6313] = 8'd105;
vmem[6314] = 8'd109;
vmem[6315] = 8'd101;
vmem[6316] = 8'd110;
vmem[6317] = 8'd116;
vmem[6318] = 8'd117;
vmem[6319] = 8'd109;
vmem[6320] = 8'd32;
vmem[6321] = 8'd110;
vmem[6322] = 8'd101;
vmem[6323] = 8'd99;
vmem[6324] = 8'd44;
vmem[6325] = 8'd32;
vmem[6326] = 8'd108;
vmem[6327] = 8'd111;
vmem[6328] = 8'd98;
vmem[6329] = 8'd111;
vmem[6330] = 8'd114;
vmem[6331] = 8'd116;
vmem[6332] = 8'd105;
vmem[6333] = 8'd115;
vmem[6334] = 8'd32;
vmem[6335] = 8'd118;
vmem[6336] = 8'd105;
vmem[6337] = 8'd116;
vmem[6338] = 8'd97;
vmem[6339] = 8'd101;
vmem[6340] = 8'd32;
vmem[6341] = 8'd101;
vmem[6342] = 8'd108;
vmem[6343] = 8'd105;
vmem[6344] = 8'd116;
vmem[6345] = 8'd46;
vmem[6346] = 8'd32;
vmem[6347] = 8'd70;
vmem[6348] = 8'd117;
vmem[6349] = 8'd115;
vmem[6350] = 8'd99;
vmem[6351] = 8'd101;
vmem[6352] = 8'd32;
vmem[6353] = 8'd117;
vmem[6354] = 8'd116;
vmem[6355] = 8'd32;
vmem[6356] = 8'd109;
vmem[6357] = 8'd97;
vmem[6358] = 8'd117;
vmem[6359] = 8'd114;
vmem[6360] = 8'd105;
vmem[6361] = 8'd115;
vmem[6362] = 8'd32;
vmem[6363] = 8'd113;
vmem[6364] = 8'd117;
vmem[6365] = 8'd105;
vmem[6366] = 8'd115;
vmem[6367] = 8'd32;
vmem[6368] = 8'd109;
vmem[6369] = 8'd101;
vmem[6370] = 8'd116;
vmem[6371] = 8'd117;
vmem[6372] = 8'd115;
vmem[6373] = 8'd32;
vmem[6374] = 8'd114;
vmem[6375] = 8'd117;
vmem[6376] = 8'd116;
vmem[6377] = 8'd114;
vmem[6378] = 8'd117;
vmem[6379] = 8'd109;
vmem[6380] = 8'd32;
vmem[6381] = 8'd102;
vmem[6382] = 8'd97;
vmem[6383] = 8'd117;
vmem[6384] = 8'd99;
vmem[6385] = 8'd105;
vmem[6386] = 8'd98;
vmem[6387] = 8'd117;
vmem[6388] = 8'd115;
vmem[6389] = 8'd46;
vmem[6390] = 8'd32;
vmem[6391] = 8'd78;
vmem[6392] = 8'd117;
vmem[6393] = 8'd108;
vmem[6394] = 8'd108;
vmem[6395] = 8'd97;
vmem[6396] = 8'd32;
vmem[6397] = 8'd108;
vmem[6398] = 8'd117;
vmem[6399] = 8'd99;
vmem[6400] = 8'd116;
vmem[6401] = 8'd117;
vmem[6402] = 8'd115;
vmem[6403] = 8'd32;
vmem[6404] = 8'd97;
vmem[6405] = 8'd114;
vmem[6406] = 8'd99;
vmem[6407] = 8'd117;
vmem[6408] = 8'd32;
vmem[6409] = 8'd105;
vmem[6410] = 8'd110;
vmem[6411] = 8'd32;
vmem[6412] = 8'd108;
vmem[6413] = 8'd111;
vmem[6414] = 8'd114;
vmem[6415] = 8'd101;
vmem[6416] = 8'd109;
vmem[6417] = 8'd32;
vmem[6418] = 8'd109;
vmem[6419] = 8'd97;
vmem[6420] = 8'd116;
vmem[6421] = 8'd116;
vmem[6422] = 8'd105;
vmem[6423] = 8'd115;
vmem[6424] = 8'd32;
vmem[6425] = 8'd117;
vmem[6426] = 8'd108;
vmem[6427] = 8'd108;
vmem[6428] = 8'd97;
vmem[6429] = 8'd109;
vmem[6430] = 8'd99;
vmem[6431] = 8'd111;
vmem[6432] = 8'd114;
vmem[6433] = 8'd112;
vmem[6434] = 8'd101;
vmem[6435] = 8'd114;
vmem[6436] = 8'd46;
vmem[6437] = 8'd32;
vmem[6438] = 8'd68;
vmem[6439] = 8'd111;
vmem[6440] = 8'd110;
vmem[6441] = 8'd101;
vmem[6442] = 8'd99;
vmem[6443] = 8'd32;
vmem[6444] = 8'd118;
vmem[6445] = 8'd105;
vmem[6446] = 8'd116;
vmem[6447] = 8'd97;
vmem[6448] = 8'd101;
vmem[6449] = 8'd32;
vmem[6450] = 8'd112;
vmem[6451] = 8'd117;
vmem[6452] = 8'd114;
vmem[6453] = 8'd117;
vmem[6454] = 8'd115;
vmem[6455] = 8'd32;
vmem[6456] = 8'd109;
vmem[6457] = 8'd101;
vmem[6458] = 8'd116;
vmem[6459] = 8'd117;
vmem[6460] = 8'd115;
vmem[6461] = 8'd46;
vmem[6462] = 8'd32;
vmem[6463] = 8'd83;
vmem[6464] = 8'd101;
vmem[6465] = 8'd100;
vmem[6466] = 8'd32;
vmem[6467] = 8'd101;
vmem[6468] = 8'd103;
vmem[6469] = 8'd101;
vmem[6470] = 8'd115;
vmem[6471] = 8'd116;
vmem[6472] = 8'd97;
vmem[6473] = 8'd115;
vmem[6474] = 8'd32;
vmem[6475] = 8'd115;
vmem[6476] = 8'd97;
vmem[6477] = 8'd112;
vmem[6478] = 8'd105;
vmem[6479] = 8'd101;
vmem[6480] = 8'd110;
vmem[6481] = 8'd32;
vmem[6482] = 8'd99;
vmem[6483] = 8'd117;
vmem[6484] = 8'd114;
vmem[6485] = 8'd115;
vmem[6486] = 8'd117;
vmem[6487] = 8'd115;
vmem[6488] = 8'd32;
vmem[6489] = 8'd108;
vmem[6490] = 8'd105;
vmem[6491] = 8'd103;
vmem[6492] = 8'd117;
vmem[6493] = 8'd108;
vmem[6494] = 8'd97;
vmem[6495] = 8'd32;
vmem[6496] = 8'd118;
vmem[6497] = 8'd101;
vmem[6498] = 8'd110;
vmem[6499] = 8'd101;
vmem[6500] = 8'd110;
vmem[6501] = 8'd97;
vmem[6502] = 8'd116;
vmem[6503] = 8'd105;
vmem[6504] = 8'd115;
vmem[6505] = 8'd32;
vmem[6506] = 8'd109;
vmem[6507] = 8'd97;
vmem[6508] = 8'd120;
vmem[6509] = 8'd105;
vmem[6510] = 8'd109;
vmem[6511] = 8'd117;
vmem[6512] = 8'd115;
vmem[6513] = 8'd46;
vmem[6514] = 8'd32;
vmem[6515] = 8'd86;
vmem[6516] = 8'd101;
vmem[6517] = 8'd115;
vmem[6518] = 8'd116;
vmem[6519] = 8'd105;
vmem[6520] = 8'd98;
vmem[6521] = 8'd117;
vmem[6522] = 8'd108;
vmem[6523] = 8'd117;
vmem[6524] = 8'd109;
vmem[6525] = 8'd32;
vmem[6526] = 8'd118;
vmem[6527] = 8'd101;
vmem[6528] = 8'd108;
vmem[6529] = 8'd32;
vmem[6530] = 8'd101;
vmem[6531] = 8'd108;
vmem[6532] = 8'd101;
vmem[6533] = 8'd105;
vmem[6534] = 8'd102;
vmem[6535] = 8'd101;
vmem[6536] = 8'd110;
vmem[6537] = 8'd100;
vmem[6538] = 8'd32;
vmem[6539] = 8'd110;
vmem[6540] = 8'd117;
vmem[6541] = 8'd110;
vmem[6542] = 8'd99;
vmem[6543] = 8'd44;
vmem[6544] = 8'd32;
vmem[6545] = 8'd115;
vmem[6546] = 8'd105;
vmem[6547] = 8'd116;
vmem[6548] = 8'd32;
vmem[6549] = 8'd97;
vmem[6550] = 8'd109;
vmem[6551] = 8'd101;
vmem[6552] = 8'd116;
vmem[6553] = 8'd32;
vmem[6554] = 8'd112;
vmem[6555] = 8'd114;
vmem[6556] = 8'd101;
vmem[6557] = 8'd116;
vmem[6558] = 8'd105;
vmem[6559] = 8'd117;
vmem[6560] = 8'd109;
vmem[6561] = 8'd32;
vmem[6562] = 8'd110;
vmem[6563] = 8'd105;
vmem[6564] = 8'd98;
vmem[6565] = 8'd104;
vmem[6566] = 8'd46;
vmem[6567] = 8'd32;
vmem[6568] = 8'd73;
vmem[6569] = 8'd110;
vmem[6570] = 8'd32;
vmem[6571] = 8'd104;
vmem[6572] = 8'd97;
vmem[6573] = 8'd99;
vmem[6574] = 8'd32;
vmem[6575] = 8'd104;
vmem[6576] = 8'd97;
vmem[6577] = 8'd98;
vmem[6578] = 8'd105;
vmem[6579] = 8'd116;
vmem[6580] = 8'd97;
vmem[6581] = 8'd115;
vmem[6582] = 8'd115;
vmem[6583] = 8'd101;
vmem[6584] = 8'd32;
vmem[6585] = 8'd112;
vmem[6586] = 8'd108;
vmem[6587] = 8'd97;
vmem[6588] = 8'd116;
vmem[6589] = 8'd101;
vmem[6590] = 8'd97;
vmem[6591] = 8'd32;
vmem[6592] = 8'd100;
vmem[6593] = 8'd105;
vmem[6594] = 8'd99;
vmem[6595] = 8'd116;
vmem[6596] = 8'd117;
vmem[6597] = 8'd109;
vmem[6598] = 8'd115;
vmem[6599] = 8'd116;
vmem[6600] = 8'd46;
vmem[6601] = 8'd32;
vmem[6602] = 8'd83;
vmem[6603] = 8'd101;
vmem[6604] = 8'd100;
vmem[6605] = 8'd32;
vmem[6606] = 8'd108;
vmem[6607] = 8'd101;
vmem[6608] = 8'd99;
vmem[6609] = 8'd116;
vmem[6610] = 8'd117;
vmem[6611] = 8'd115;
vmem[6612] = 8'd32;
vmem[6613] = 8'd97;
vmem[6614] = 8'd110;
vmem[6615] = 8'd116;
vmem[6616] = 8'd101;
vmem[6617] = 8'd44;
vmem[6618] = 8'd32;
vmem[6619] = 8'd102;
vmem[6620] = 8'd114;
vmem[6621] = 8'd105;
vmem[6622] = 8'd110;
vmem[6623] = 8'd103;
vmem[6624] = 8'd105;
vmem[6625] = 8'd108;
vmem[6626] = 8'd108;
vmem[6627] = 8'd97;
vmem[6628] = 8'd32;
vmem[6629] = 8'd118;
vmem[6630] = 8'd101;
vmem[6631] = 8'd108;
vmem[6632] = 8'd32;
vmem[6633] = 8'd100;
vmem[6634] = 8'd111;
vmem[6635] = 8'd108;
vmem[6636] = 8'd111;
vmem[6637] = 8'd114;
vmem[6638] = 8'd32;
vmem[6639] = 8'd118;
vmem[6640] = 8'd105;
vmem[6641] = 8'd116;
vmem[6642] = 8'd97;
vmem[6643] = 8'd101;
vmem[6644] = 8'd44;
vmem[6645] = 8'd32;
vmem[6646] = 8'd116;
vmem[6647] = 8'd101;
vmem[6648] = 8'd109;
vmem[6649] = 8'd112;
vmem[6650] = 8'd111;
vmem[6651] = 8'd114;
vmem[6652] = 8'd32;
vmem[6653] = 8'd99;
vmem[6654] = 8'd111;
vmem[6655] = 8'd109;
vmem[6656] = 8'd109;
vmem[6657] = 8'd111;
vmem[6658] = 8'd100;
vmem[6659] = 8'd111;
vmem[6660] = 8'd32;
vmem[6661] = 8'd108;
vmem[6662] = 8'd97;
vmem[6663] = 8'd99;
vmem[6664] = 8'd117;
vmem[6665] = 8'd115;
vmem[6666] = 8'd46;
vmem[6667] = 8'd32;
vmem[6668] = 8'd77;
vmem[6669] = 8'd111;
vmem[6670] = 8'd114;
vmem[6671] = 8'd98;
vmem[6672] = 8'd105;
vmem[6673] = 8'd32;
vmem[6674] = 8'd97;
vmem[6675] = 8'd99;
vmem[6676] = 8'd99;
vmem[6677] = 8'd117;
vmem[6678] = 8'd109;
vmem[6679] = 8'd115;
vmem[6680] = 8'd97;
vmem[6681] = 8'd110;
vmem[6682] = 8'd44;
vmem[6683] = 8'd32;
vmem[6684] = 8'd116;
vmem[6685] = 8'd101;
vmem[6686] = 8'd108;
vmem[6687] = 8'd108;
vmem[6688] = 8'd117;
vmem[6689] = 8'd115;
vmem[6690] = 8'd32;
vmem[6691] = 8'd100;
vmem[6692] = 8'd105;
vmem[6693] = 8'd99;
vmem[6694] = 8'd116;
vmem[6695] = 8'd117;
vmem[6696] = 8'd109;
vmem[6697] = 8'd32;
vmem[6698] = 8'd102;
vmem[6699] = 8'd114;
vmem[6700] = 8'd105;
vmem[6701] = 8'd110;
vmem[6702] = 8'd103;
vmem[6703] = 8'd105;
vmem[6704] = 8'd108;
vmem[6705] = 8'd108;
vmem[6706] = 8'd97;
vmem[6707] = 8'd32;
vmem[6708] = 8'd115;
vmem[6709] = 8'd97;
vmem[6710] = 8'd103;
vmem[6711] = 8'd105;
vmem[6712] = 8'd116;
vmem[6713] = 8'd116;
vmem[6714] = 8'd105;
vmem[6715] = 8'd115;
vmem[6716] = 8'd44;
vmem[6717] = 8'd32;
vmem[6718] = 8'd111;
vmem[6719] = 8'd100;
vmem[6720] = 8'd105;
vmem[6721] = 8'd111;
vmem[6722] = 8'd32;
vmem[6723] = 8'd97;
vmem[6724] = 8'd110;
vmem[6725] = 8'd116;
vmem[6726] = 8'd101;
vmem[6727] = 8'd32;
vmem[6728] = 8'd109;
vmem[6729] = 8'd97;
vmem[6730] = 8'd108;
vmem[6731] = 8'd101;
vmem[6732] = 8'd115;
vmem[6733] = 8'd117;
vmem[6734] = 8'd97;
vmem[6735] = 8'd100;
vmem[6736] = 8'd97;
vmem[6737] = 8'd32;
vmem[6738] = 8'd117;
vmem[6739] = 8'd114;
vmem[6740] = 8'd110;
vmem[6741] = 8'd97;
vmem[6742] = 8'd44;
vmem[6743] = 8'd32;
vmem[6744] = 8'd110;
vmem[6745] = 8'd101;
vmem[6746] = 8'd99;
vmem[6747] = 8'd32;
vmem[6748] = 8'd101;
vmem[6749] = 8'd108;
vmem[6750] = 8'd101;
vmem[6751] = 8'd109;
vmem[6752] = 8'd101;
vmem[6753] = 8'd110;
vmem[6754] = 8'd116;
vmem[6755] = 8'd117;
vmem[6756] = 8'd109;
vmem[6757] = 8'd32;
vmem[6758] = 8'd116;
vmem[6759] = 8'd117;
vmem[6760] = 8'd114;
vmem[6761] = 8'd112;
vmem[6762] = 8'd105;
vmem[6763] = 8'd115;
vmem[6764] = 8'd32;
vmem[6765] = 8'd109;
vmem[6766] = 8'd97;
vmem[6767] = 8'd103;
vmem[6768] = 8'd110;
vmem[6769] = 8'd97;
vmem[6770] = 8'd32;
vmem[6771] = 8'd97;
vmem[6772] = 8'd32;
vmem[6773] = 8'd105;
vmem[6774] = 8'd112;
vmem[6775] = 8'd115;
vmem[6776] = 8'd117;
vmem[6777] = 8'd109;
vmem[6778] = 8'd46;
vmem[6779] = 8'd32;
vmem[6780] = 8'd68;
vmem[6781] = 8'd117;
vmem[6782] = 8'd105;
vmem[6783] = 8'd115;
vmem[6784] = 8'd32;
vmem[6785] = 8'd115;
vmem[6786] = 8'd101;
vmem[6787] = 8'd100;
vmem[6788] = 8'd32;
vmem[6789] = 8'd97;
vmem[6790] = 8'd117;
vmem[6791] = 8'd103;
vmem[6792] = 8'd117;
vmem[6793] = 8'd101;
vmem[6794] = 8'd32;
vmem[6795] = 8'd101;
vmem[6796] = 8'd108;
vmem[6797] = 8'd105;
vmem[6798] = 8'd116;
vmem[6799] = 8'd46;
vmem[6800] = 8'd32;
vmem[6801] = 8'd67;
vmem[6802] = 8'd114;
vmem[6803] = 8'd97;
vmem[6804] = 8'd115;
vmem[6805] = 8'd32;
vmem[6806] = 8'd117;
vmem[6807] = 8'd108;
vmem[6808] = 8'd116;
vmem[6809] = 8'd114;
vmem[6810] = 8'd105;
vmem[6811] = 8'd99;
vmem[6812] = 8'd105;
vmem[6813] = 8'd101;
vmem[6814] = 8'd115;
vmem[6815] = 8'd32;
vmem[6816] = 8'd101;
vmem[6817] = 8'd115;
vmem[6818] = 8'd116;
vmem[6819] = 8'd32;
vmem[6820] = 8'd101;
vmem[6821] = 8'd116;
vmem[6822] = 8'd32;
vmem[6823] = 8'd97;
vmem[6824] = 8'd114;
vmem[6825] = 8'd99;
vmem[6826] = 8'd117;
vmem[6827] = 8'd32;
vmem[6828] = 8'd112;
vmem[6829] = 8'd117;
vmem[6830] = 8'd108;
vmem[6831] = 8'd118;
vmem[6832] = 8'd105;
vmem[6833] = 8'd110;
vmem[6834] = 8'd97;
vmem[6835] = 8'd114;
vmem[6836] = 8'd32;
vmem[6837] = 8'd112;
vmem[6838] = 8'd117;
vmem[6839] = 8'd108;
vmem[6840] = 8'd118;
vmem[6841] = 8'd105;
vmem[6842] = 8'd110;
vmem[6843] = 8'd97;
vmem[6844] = 8'd114;
vmem[6845] = 8'd46;
vmem[6846] = 8'd32;
vmem[6847] = 8'd67;
vmem[6848] = 8'd117;
vmem[6849] = 8'd114;
vmem[6850] = 8'd97;
vmem[6851] = 8'd98;
vmem[6852] = 8'd105;
vmem[6853] = 8'd116;
vmem[6854] = 8'd117;
vmem[6855] = 8'd114;
vmem[6856] = 8'd32;
vmem[6857] = 8'd109;
vmem[6858] = 8'd97;
vmem[6859] = 8'd117;
vmem[6860] = 8'd114;
vmem[6861] = 8'd105;
vmem[6862] = 8'd115;
vmem[6863] = 8'd32;
vmem[6864] = 8'd109;
vmem[6865] = 8'd97;
vmem[6866] = 8'd115;
vmem[6867] = 8'd115;
vmem[6868] = 8'd97;
vmem[6869] = 8'd44;
vmem[6870] = 8'd32;
vmem[6871] = 8'd115;
vmem[6872] = 8'd97;
vmem[6873] = 8'd103;
vmem[6874] = 8'd105;
vmem[6875] = 8'd116;
vmem[6876] = 8'd116;
vmem[6877] = 8'd105;
vmem[6878] = 8'd115;
vmem[6879] = 8'd32;
vmem[6880] = 8'd118;
vmem[6881] = 8'd101;
vmem[6882] = 8'd108;
vmem[6883] = 8'd32;
vmem[6884] = 8'd109;
vmem[6885] = 8'd111;
vmem[6886] = 8'd108;
vmem[6887] = 8'd108;
vmem[6888] = 8'd105;
vmem[6889] = 8'd115;
vmem[6890] = 8'd32;
vmem[6891] = 8'd113;
vmem[6892] = 8'd117;
vmem[6893] = 8'd105;
vmem[6894] = 8'd115;
vmem[6895] = 8'd44;
vmem[6896] = 8'd32;
vmem[6897] = 8'd109;
vmem[6898] = 8'd97;
vmem[6899] = 8'd108;
vmem[6900] = 8'd101;
vmem[6901] = 8'd115;
vmem[6902] = 8'd117;
vmem[6903] = 8'd97;
vmem[6904] = 8'd100;
vmem[6905] = 8'd97;
vmem[6906] = 8'd32;
vmem[6907] = 8'd110;
vmem[6908] = 8'd101;
vmem[6909] = 8'd99;
vmem[6910] = 8'd32;
vmem[6911] = 8'd116;
vmem[6912] = 8'd111;
vmem[6913] = 8'd114;
vmem[6914] = 8'd116;
vmem[6915] = 8'd111;
vmem[6916] = 8'd114;
vmem[6917] = 8'd46;
vmem[6918] = 8'd32;
vmem[6919] = 8'd65;
vmem[6920] = 8'd108;
vmem[6921] = 8'd105;
vmem[6922] = 8'd113;
vmem[6923] = 8'd117;
vmem[6924] = 8'd97;
vmem[6925] = 8'd109;
vmem[6926] = 8'd32;
vmem[6927] = 8'd102;
vmem[6928] = 8'd97;
vmem[6929] = 8'd117;
vmem[6930] = 8'd99;
vmem[6931] = 8'd105;
vmem[6932] = 8'd98;
vmem[6933] = 8'd117;
vmem[6934] = 8'd115;
vmem[6935] = 8'd32;
vmem[6936] = 8'd117;
vmem[6937] = 8'd116;
vmem[6938] = 8'd32;
vmem[6939] = 8'd113;
vmem[6940] = 8'd117;
vmem[6941] = 8'd97;
vmem[6942] = 8'd109;
vmem[6943] = 8'd32;
vmem[6944] = 8'd110;
vmem[6945] = 8'd111;
vmem[6946] = 8'd110;
vmem[6947] = 8'd32;
vmem[6948] = 8'd104;
vmem[6949] = 8'd101;
vmem[6950] = 8'd110;
vmem[6951] = 8'd100;
vmem[6952] = 8'd114;
vmem[6953] = 8'd101;
vmem[6954] = 8'd114;
vmem[6955] = 8'd105;
vmem[6956] = 8'd116;
vmem[6957] = 8'd46;
vmem[6958] = 8'd32;
vmem[6959] = 8'd77;
vmem[6960] = 8'd111;
vmem[6961] = 8'd114;
vmem[6962] = 8'd98;
vmem[6963] = 8'd105;
vmem[6964] = 8'd32;
vmem[6965] = 8'd118;
vmem[6966] = 8'd101;
vmem[6967] = 8'd104;
vmem[6968] = 8'd105;
vmem[6969] = 8'd99;
vmem[6970] = 8'd117;
vmem[6971] = 8'd108;
vmem[6972] = 8'd97;
vmem[6973] = 8'd32;
vmem[6974] = 8'd99;
vmem[6975] = 8'd111;
vmem[6976] = 8'd109;
vmem[6977] = 8'd109;
vmem[6978] = 8'd111;
vmem[6979] = 8'd100;
vmem[6980] = 8'd111;
vmem[6981] = 8'd32;
vmem[6982] = 8'd108;
vmem[6983] = 8'd105;
vmem[6984] = 8'd98;
vmem[6985] = 8'd101;
vmem[6986] = 8'd114;
vmem[6987] = 8'd111;
vmem[6988] = 8'd46;
vmem[6989] = 8'd32;
vmem[6990] = 8'd67;
vmem[6991] = 8'd117;
vmem[6992] = 8'd114;
vmem[6993] = 8'd97;
vmem[6994] = 8'd98;
vmem[6995] = 8'd105;
vmem[6996] = 8'd116;
vmem[6997] = 8'd117;
vmem[6998] = 8'd114;
vmem[6999] = 8'd32;
vmem[7000] = 8'd115;
vmem[7001] = 8'd105;
vmem[7002] = 8'd116;
vmem[7003] = 8'd32;
vmem[7004] = 8'd97;
vmem[7005] = 8'd109;
vmem[7006] = 8'd101;
vmem[7007] = 8'd116;
vmem[7008] = 8'd32;
vmem[7009] = 8'd102;
vmem[7010] = 8'd105;
vmem[7011] = 8'd110;
vmem[7012] = 8'd105;
vmem[7013] = 8'd98;
vmem[7014] = 8'd117;
vmem[7015] = 8'd115;
vmem[7016] = 8'd32;
vmem[7017] = 8'd116;
vmem[7018] = 8'd101;
vmem[7019] = 8'd108;
vmem[7020] = 8'd108;
vmem[7021] = 8'd117;
vmem[7022] = 8'd115;
vmem[7023] = 8'd46;
vmem[7024] = 8'd32;
vmem[7025] = 8'd83;
vmem[7026] = 8'd101;
vmem[7027] = 8'd100;
vmem[7028] = 8'd32;
vmem[7029] = 8'd110;
vmem[7030] = 8'd105;
vmem[7031] = 8'd115;
vmem[7032] = 8'd105;
vmem[7033] = 8'd32;
vmem[7034] = 8'd101;
vmem[7035] = 8'd114;
vmem[7036] = 8'd97;
vmem[7037] = 8'd116;
vmem[7038] = 8'd44;
vmem[7039] = 8'd32;
vmem[7040] = 8'd116;
vmem[7041] = 8'd105;
vmem[7042] = 8'd110;
vmem[7043] = 8'd99;
vmem[7044] = 8'd105;
vmem[7045] = 8'd100;
vmem[7046] = 8'd117;
vmem[7047] = 8'd110;
vmem[7048] = 8'd116;
vmem[7049] = 8'd32;
vmem[7050] = 8'd117;
vmem[7051] = 8'd116;
vmem[7052] = 8'd32;
vmem[7053] = 8'd108;
vmem[7054] = 8'd97;
vmem[7055] = 8'd111;
vmem[7056] = 8'd114;
vmem[7057] = 8'd101;
vmem[7058] = 8'd101;
vmem[7059] = 8'd116;
vmem[7060] = 8'd32;
vmem[7061] = 8'd115;
vmem[7062] = 8'd105;
vmem[7063] = 8'd116;
vmem[7064] = 8'd32;
vmem[7065] = 8'd97;
vmem[7066] = 8'd109;
vmem[7067] = 8'd101;
vmem[7068] = 8'd116;
vmem[7069] = 8'd44;
vmem[7070] = 8'd32;
vmem[7071] = 8'd101;
vmem[7072] = 8'd108;
vmem[7073] = 8'd101;
vmem[7074] = 8'd109;
vmem[7075] = 8'd101;
vmem[7076] = 8'd110;
vmem[7077] = 8'd116;
vmem[7078] = 8'd117;
vmem[7079] = 8'd109;
vmem[7080] = 8'd32;
vmem[7081] = 8'd118;
vmem[7082] = 8'd101;
vmem[7083] = 8'd108;
vmem[7084] = 8'd32;
vmem[7085] = 8'd108;
vmem[7086] = 8'd111;
vmem[7087] = 8'd114;
vmem[7088] = 8'd101;
vmem[7089] = 8'd109;
vmem[7090] = 8'd46;
vmem[7091] = 8'd32;
vmem[7092] = 8'd68;
vmem[7093] = 8'd111;
vmem[7094] = 8'd110;
vmem[7095] = 8'd101;
vmem[7096] = 8'd99;
vmem[7097] = 8'd32;
vmem[7098] = 8'd97;
vmem[7099] = 8'd116;
vmem[7100] = 8'd32;
vmem[7101] = 8'd110;
vmem[7102] = 8'd117;
vmem[7103] = 8'd110;
vmem[7104] = 8'd99;
vmem[7105] = 8'd32;
vmem[7106] = 8'd110;
vmem[7107] = 8'd101;
vmem[7108] = 8'd99;
vmem[7109] = 8'd32;
vmem[7110] = 8'd108;
vmem[7111] = 8'd105;
vmem[7112] = 8'd98;
vmem[7113] = 8'd101;
vmem[7114] = 8'd114;
vmem[7115] = 8'd111;
vmem[7116] = 8'd32;
vmem[7117] = 8'd116;
vmem[7118] = 8'd101;
vmem[7119] = 8'd109;
vmem[7120] = 8'd112;
vmem[7121] = 8'd117;
vmem[7122] = 8'd115;
vmem[7123] = 8'd32;
vmem[7124] = 8'd115;
vmem[7125] = 8'd101;
vmem[7126] = 8'd109;
vmem[7127] = 8'd112;
vmem[7128] = 8'd101;
vmem[7129] = 8'd114;
vmem[7130] = 8'd32;
vmem[7131] = 8'd117;
vmem[7132] = 8'd116;
vmem[7133] = 8'd32;
vmem[7134] = 8'd105;
vmem[7135] = 8'd100;
vmem[7136] = 8'd32;
vmem[7137] = 8'd100;
vmem[7138] = 8'd105;
vmem[7139] = 8'd97;
vmem[7140] = 8'd109;
vmem[7141] = 8'd46;
vmem[7142] = 8'd32;
vmem[7143] = 8'd65;
vmem[7144] = 8'd101;
vmem[7145] = 8'd110;
vmem[7146] = 8'd101;
vmem[7147] = 8'd97;
vmem[7148] = 8'd110;
vmem[7149] = 8'd32;
vmem[7150] = 8'd99;
vmem[7151] = 8'd111;
vmem[7152] = 8'd109;
vmem[7153] = 8'd109;
vmem[7154] = 8'd111;
vmem[7155] = 8'd100;
vmem[7156] = 8'd111;
vmem[7157] = 8'd32;
vmem[7158] = 8'd98;
vmem[7159] = 8'd108;
vmem[7160] = 8'd97;
vmem[7161] = 8'd110;
vmem[7162] = 8'd100;
vmem[7163] = 8'd105;
vmem[7164] = 8'd116;
vmem[7165] = 8'd32;
vmem[7166] = 8'd101;
vmem[7167] = 8'd110;
vmem[7168] = 8'd105;
vmem[7169] = 8'd109;
vmem[7170] = 8'd44;
vmem[7171] = 8'd32;
vmem[7172] = 8'd115;
vmem[7173] = 8'd101;
vmem[7174] = 8'd100;
vmem[7175] = 8'd32;
vmem[7176] = 8'd104;
vmem[7177] = 8'd101;
vmem[7178] = 8'd110;
vmem[7179] = 8'd100;
vmem[7180] = 8'd114;
vmem[7181] = 8'd101;
vmem[7182] = 8'd114;
vmem[7183] = 8'd105;
vmem[7184] = 8'd116;
vmem[7185] = 8'd32;
vmem[7186] = 8'd105;
vmem[7187] = 8'd112;
vmem[7188] = 8'd115;
vmem[7189] = 8'd117;
vmem[7190] = 8'd109;
vmem[7191] = 8'd32;
vmem[7192] = 8'd102;
vmem[7193] = 8'd101;
vmem[7194] = 8'd114;
vmem[7195] = 8'd109;
vmem[7196] = 8'd101;
vmem[7197] = 8'd110;
vmem[7198] = 8'd116;
vmem[7199] = 8'd117;
vmem[7200] = 8'd109;
vmem[7201] = 8'd32;
vmem[7202] = 8'd115;
vmem[7203] = 8'd101;
vmem[7204] = 8'd100;
vmem[7205] = 8'd46;
vmem[7206] = 8'd32;
vmem[7207] = 8'd70;
vmem[7208] = 8'd117;
vmem[7209] = 8'd115;
vmem[7210] = 8'd99;
vmem[7211] = 8'd101;
vmem[7212] = 8'd32;
vmem[7213] = 8'd97;
vmem[7214] = 8'd32;
vmem[7215] = 8'd109;
vmem[7216] = 8'd101;
vmem[7217] = 8'd116;
vmem[7218] = 8'd117;
vmem[7219] = 8'd115;
vmem[7220] = 8'd32;
vmem[7221] = 8'd110;
vmem[7222] = 8'd101;
vmem[7223] = 8'd99;
vmem[7224] = 8'd32;
vmem[7225] = 8'd110;
vmem[7226] = 8'd105;
vmem[7227] = 8'd115;
vmem[7228] = 8'd108;
vmem[7229] = 8'd32;
vmem[7230] = 8'd101;
vmem[7231] = 8'd102;
vmem[7232] = 8'd102;
vmem[7233] = 8'd105;
vmem[7234] = 8'd99;
vmem[7235] = 8'd105;
vmem[7236] = 8'd116;
vmem[7237] = 8'd117;
vmem[7238] = 8'd114;
vmem[7239] = 8'd32;
vmem[7240] = 8'd108;
vmem[7241] = 8'd117;
vmem[7242] = 8'd99;
vmem[7243] = 8'd116;
vmem[7244] = 8'd117;
vmem[7245] = 8'd115;
vmem[7246] = 8'd32;
vmem[7247] = 8'd97;
vmem[7248] = 8'd116;
vmem[7249] = 8'd32;
vmem[7250] = 8'd97;
vmem[7251] = 8'd116;
vmem[7252] = 8'd32;
vmem[7253] = 8'd108;
vmem[7254] = 8'd97;
vmem[7255] = 8'd99;
vmem[7256] = 8'd117;
vmem[7257] = 8'd115;
vmem[7258] = 8'd46;
vmem[7259] = 8'd32;
vmem[7260] = 8'd77;
vmem[7261] = 8'd97;
vmem[7262] = 8'd117;
vmem[7263] = 8'd114;
vmem[7264] = 8'd105;
vmem[7265] = 8'd115;
vmem[7266] = 8'd32;
vmem[7267] = 8'd108;
vmem[7268] = 8'd97;
vmem[7269] = 8'd99;
vmem[7270] = 8'd105;
vmem[7271] = 8'd110;
vmem[7272] = 8'd105;
vmem[7273] = 8'd97;
vmem[7274] = 8'd32;
vmem[7275] = 8'd110;
vmem[7276] = 8'd105;
vmem[7277] = 8'd115;
vmem[7278] = 8'd108;
vmem[7279] = 8'd32;
vmem[7280] = 8'd100;
vmem[7281] = 8'd105;
vmem[7282] = 8'd97;
vmem[7283] = 8'd109;
vmem[7284] = 8'd44;
vmem[7285] = 8'd32;
vmem[7286] = 8'd101;
vmem[7287] = 8'd103;
vmem[7288] = 8'd101;
vmem[7289] = 8'd116;
vmem[7290] = 8'd32;
vmem[7291] = 8'd116;
vmem[7292] = 8'd114;
vmem[7293] = 8'd105;
vmem[7294] = 8'd115;
vmem[7295] = 8'd116;
vmem[7296] = 8'd105;
vmem[7297] = 8'd113;
vmem[7298] = 8'd117;
vmem[7299] = 8'd101;
vmem[7300] = 8'd32;
vmem[7301] = 8'd108;
vmem[7302] = 8'd97;
vmem[7303] = 8'd99;
vmem[7304] = 8'd117;
vmem[7305] = 8'd115;
vmem[7306] = 8'd32;
vmem[7307] = 8'd99;
vmem[7308] = 8'd111;
vmem[7309] = 8'd110;
vmem[7310] = 8'd115;
vmem[7311] = 8'd101;
vmem[7312] = 8'd113;
vmem[7313] = 8'd117;
vmem[7314] = 8'd97;
vmem[7315] = 8'd116;
vmem[7316] = 8'd32;
vmem[7317] = 8'd115;
vmem[7318] = 8'd105;
vmem[7319] = 8'd116;
vmem[7320] = 8'd32;
vmem[7321] = 8'd97;
vmem[7322] = 8'd109;
vmem[7323] = 8'd101;
vmem[7324] = 8'd116;
vmem[7325] = 8'd46;
vmem[7326] = 8'd32;
vmem[7327] = 8'd80;
vmem[7328] = 8'd114;
vmem[7329] = 8'd97;
vmem[7330] = 8'd101;
vmem[7331] = 8'd115;
vmem[7332] = 8'd101;
vmem[7333] = 8'd110;
vmem[7334] = 8'd116;
vmem[7335] = 8'd32;
vmem[7336] = 8'd117;
vmem[7337] = 8'd108;
vmem[7338] = 8'd108;
vmem[7339] = 8'd97;
vmem[7340] = 8'd109;
vmem[7341] = 8'd99;
vmem[7342] = 8'd111;
vmem[7343] = 8'd114;
vmem[7344] = 8'd112;
vmem[7345] = 8'd101;
vmem[7346] = 8'd114;
vmem[7347] = 8'd32;
vmem[7348] = 8'd102;
vmem[7349] = 8'd101;
vmem[7350] = 8'd108;
vmem[7351] = 8'd105;
vmem[7352] = 8'd115;
vmem[7353] = 8'd32;
vmem[7354] = 8'd115;
vmem[7355] = 8'd101;
vmem[7356] = 8'd100;
vmem[7357] = 8'd32;
vmem[7358] = 8'd113;
vmem[7359] = 8'd117;
vmem[7360] = 8'd97;
vmem[7361] = 8'd109;
vmem[7362] = 8'd32;
vmem[7363] = 8'd112;
vmem[7364] = 8'd117;
vmem[7365] = 8'd108;
vmem[7366] = 8'd118;
vmem[7367] = 8'd105;
vmem[7368] = 8'd110;
vmem[7369] = 8'd97;
vmem[7370] = 8'd114;
vmem[7371] = 8'd32;
vmem[7372] = 8'd116;
vmem[7373] = 8'd114;
vmem[7374] = 8'd105;
vmem[7375] = 8'd115;
vmem[7376] = 8'd116;
vmem[7377] = 8'd105;
vmem[7378] = 8'd113;
vmem[7379] = 8'd117;
vmem[7380] = 8'd101;
vmem[7381] = 8'd46;
vmem[7382] = 8'd32;
vmem[7383] = 8'd78;
vmem[7384] = 8'd117;
vmem[7385] = 8'd108;
vmem[7386] = 8'd108;
vmem[7387] = 8'd97;
vmem[7388] = 8'd109;
vmem[7389] = 8'd32;
vmem[7390] = 8'd116;
vmem[7391] = 8'd105;
vmem[7392] = 8'd110;
vmem[7393] = 8'd99;
vmem[7394] = 8'd105;
vmem[7395] = 8'd100;
vmem[7396] = 8'd117;
vmem[7397] = 8'd110;
vmem[7398] = 8'd116;
vmem[7399] = 8'd32;
vmem[7400] = 8'd103;
vmem[7401] = 8'd114;
vmem[7402] = 8'd97;
vmem[7403] = 8'd118;
vmem[7404] = 8'd105;
vmem[7405] = 8'd100;
vmem[7406] = 8'd97;
vmem[7407] = 8'd32;
vmem[7408] = 8'd112;
vmem[7409] = 8'd117;
vmem[7410] = 8'd114;
vmem[7411] = 8'd117;
vmem[7412] = 8'd115;
vmem[7413] = 8'd32;
vmem[7414] = 8'd112;
vmem[7415] = 8'd111;
vmem[7416] = 8'd114;
vmem[7417] = 8'd116;
vmem[7418] = 8'd116;
vmem[7419] = 8'd105;
vmem[7420] = 8'd116;
vmem[7421] = 8'd111;
vmem[7422] = 8'd114;
vmem[7423] = 8'd32;
vmem[7424] = 8'd101;
vmem[7425] = 8'd117;
vmem[7426] = 8'd105;
vmem[7427] = 8'd115;
vmem[7428] = 8'd109;
vmem[7429] = 8'd111;
vmem[7430] = 8'd100;
vmem[7431] = 8'd46;
vmem[7432] = 8'd32;
vmem[7433] = 8'd86;
vmem[7434] = 8'd101;
vmem[7435] = 8'd115;
vmem[7436] = 8'd116;
vmem[7437] = 8'd105;
vmem[7438] = 8'd98;
vmem[7439] = 8'd117;
vmem[7440] = 8'd108;
vmem[7441] = 8'd117;
vmem[7442] = 8'd109;
vmem[7443] = 8'd32;
vmem[7444] = 8'd110;
vmem[7445] = 8'd101;
vmem[7446] = 8'd99;
vmem[7447] = 8'd32;
vmem[7448] = 8'd109;
vmem[7449] = 8'd101;
vmem[7450] = 8'd116;
vmem[7451] = 8'd117;
vmem[7452] = 8'd115;
vmem[7453] = 8'd32;
vmem[7454] = 8'd115;
vmem[7455] = 8'd105;
vmem[7456] = 8'd116;
vmem[7457] = 8'd32;
vmem[7458] = 8'd97;
vmem[7459] = 8'd109;
vmem[7460] = 8'd101;
vmem[7461] = 8'd116;
vmem[7462] = 8'd32;
vmem[7463] = 8'd97;
vmem[7464] = 8'd117;
vmem[7465] = 8'd103;
vmem[7466] = 8'd117;
vmem[7467] = 8'd101;
vmem[7468] = 8'd32;
vmem[7469] = 8'd115;
vmem[7470] = 8'd97;
vmem[7471] = 8'd103;
vmem[7472] = 8'd105;
vmem[7473] = 8'd116;
vmem[7474] = 8'd116;
vmem[7475] = 8'd105;
vmem[7476] = 8'd115;
vmem[7477] = 8'd32;
vmem[7478] = 8'd101;
vmem[7479] = 8'd102;
vmem[7480] = 8'd102;
vmem[7481] = 8'd105;
vmem[7482] = 8'd99;
vmem[7483] = 8'd105;
vmem[7484] = 8'd116;
vmem[7485] = 8'd117;
vmem[7486] = 8'd114;
vmem[7487] = 8'd46;
vmem[7488] = 8'd32;
vmem[7489] = 8'd80;
vmem[7490] = 8'd101;
vmem[7491] = 8'd108;
vmem[7492] = 8'd108;
vmem[7493] = 8'd101;
vmem[7494] = 8'd110;
vmem[7495] = 8'd116;
vmem[7496] = 8'd101;
vmem[7497] = 8'd115;
vmem[7498] = 8'd113;
vmem[7499] = 8'd117;
vmem[7500] = 8'd101;
vmem[7501] = 8'd32;
vmem[7502] = 8'd104;
vmem[7503] = 8'd97;
vmem[7504] = 8'd98;
vmem[7505] = 8'd105;
vmem[7506] = 8'd116;
vmem[7507] = 8'd97;
vmem[7508] = 8'd110;
vmem[7509] = 8'd116;
vmem[7510] = 8'd32;
vmem[7511] = 8'd109;
vmem[7512] = 8'd111;
vmem[7513] = 8'd114;
vmem[7514] = 8'd98;
vmem[7515] = 8'd105;
vmem[7516] = 8'd32;
vmem[7517] = 8'd116;
vmem[7518] = 8'd114;
vmem[7519] = 8'd105;
vmem[7520] = 8'd115;
vmem[7521] = 8'd116;
vmem[7522] = 8'd105;
vmem[7523] = 8'd113;
vmem[7524] = 8'd117;
vmem[7525] = 8'd101;
vmem[7526] = 8'd32;
vmem[7527] = 8'd115;
vmem[7528] = 8'd101;
vmem[7529] = 8'd110;
vmem[7530] = 8'd101;
vmem[7531] = 8'd99;
vmem[7532] = 8'd116;
vmem[7533] = 8'd117;
vmem[7534] = 8'd115;
vmem[7535] = 8'd32;
vmem[7536] = 8'd101;
vmem[7537] = 8'd116;
vmem[7538] = 8'd32;
vmem[7539] = 8'd110;
vmem[7540] = 8'd101;
vmem[7541] = 8'd116;
vmem[7542] = 8'd117;
vmem[7543] = 8'd115;
vmem[7544] = 8'd32;
vmem[7545] = 8'd101;
vmem[7546] = 8'd116;
vmem[7547] = 8'd32;
vmem[7548] = 8'd109;
vmem[7549] = 8'd97;
vmem[7550] = 8'd108;
vmem[7551] = 8'd101;
vmem[7552] = 8'd115;
vmem[7553] = 8'd117;
vmem[7554] = 8'd97;
vmem[7555] = 8'd100;
vmem[7556] = 8'd97;
vmem[7557] = 8'd32;
vmem[7558] = 8'd102;
vmem[7559] = 8'd97;
vmem[7560] = 8'd109;
vmem[7561] = 8'd101;
vmem[7562] = 8'd115;
vmem[7563] = 8'd32;
vmem[7564] = 8'd97;
vmem[7565] = 8'd99;
vmem[7566] = 8'd32;
vmem[7567] = 8'd116;
vmem[7568] = 8'd117;
vmem[7569] = 8'd114;
vmem[7570] = 8'd112;
vmem[7571] = 8'd105;
vmem[7572] = 8'd115;
vmem[7573] = 8'd32;
vmem[7574] = 8'd101;
vmem[7575] = 8'd103;
vmem[7576] = 8'd101;
vmem[7577] = 8'd115;
vmem[7578] = 8'd116;
vmem[7579] = 8'd97;
vmem[7580] = 8'd115;
vmem[7581] = 8'd46;
vmem[7582] = 8'd32;
vmem[7583] = 8'd83;
vmem[7584] = 8'd101;
vmem[7585] = 8'd100;
vmem[7586] = 8'd32;
vmem[7587] = 8'd115;
vmem[7588] = 8'd105;
vmem[7589] = 8'd116;
vmem[7590] = 8'd32;
vmem[7591] = 8'd97;
vmem[7592] = 8'd109;
vmem[7593] = 8'd101;
vmem[7594] = 8'd116;
vmem[7595] = 8'd32;
vmem[7596] = 8'd109;
vmem[7597] = 8'd101;
vmem[7598] = 8'd116;
vmem[7599] = 8'd117;
vmem[7600] = 8'd115;
vmem[7601] = 8'd32;
vmem[7602] = 8'd115;
vmem[7603] = 8'd101;
vmem[7604] = 8'd100;
vmem[7605] = 8'd32;
vmem[7606] = 8'd101;
vmem[7607] = 8'd115;
vmem[7608] = 8'd116;
vmem[7609] = 8'd32;
vmem[7610] = 8'd118;
vmem[7611] = 8'd101;
vmem[7612] = 8'd104;
vmem[7613] = 8'd105;
vmem[7614] = 8'd99;
vmem[7615] = 8'd117;
vmem[7616] = 8'd108;
vmem[7617] = 8'd97;
vmem[7618] = 8'd32;
vmem[7619] = 8'd99;
vmem[7620] = 8'd111;
vmem[7621] = 8'd110;
vmem[7622] = 8'd118;
vmem[7623] = 8'd97;
vmem[7624] = 8'd108;
vmem[7625] = 8'd108;
vmem[7626] = 8'd105;
vmem[7627] = 8'd115;
vmem[7628] = 8'd46;
vmem[7629] = 8'd32;
vmem[7630] = 8'd65;
vmem[7631] = 8'd108;
vmem[7632] = 8'd105;
vmem[7633] = 8'd113;
vmem[7634] = 8'd117;
vmem[7635] = 8'd97;
vmem[7636] = 8'd109;
vmem[7637] = 8'd32;
vmem[7638] = 8'd101;
vmem[7639] = 8'd103;
vmem[7640] = 8'd101;
vmem[7641] = 8'd116;
vmem[7642] = 8'd32;
vmem[7643] = 8'd97;
vmem[7644] = 8'd114;
vmem[7645] = 8'd99;
vmem[7646] = 8'd117;
vmem[7647] = 8'd32;
vmem[7648] = 8'd101;
vmem[7649] = 8'd108;
vmem[7650] = 8'd101;
vmem[7651] = 8'd109;
vmem[7652] = 8'd101;
vmem[7653] = 8'd110;
vmem[7654] = 8'd116;
vmem[7655] = 8'd117;
vmem[7656] = 8'd109;
vmem[7657] = 8'd44;
vmem[7658] = 8'd32;
vmem[7659] = 8'd109;
vmem[7660] = 8'd111;
vmem[7661] = 8'd108;
vmem[7662] = 8'd108;
vmem[7663] = 8'd105;
vmem[7664] = 8'd115;
vmem[7665] = 8'd32;
vmem[7666] = 8'd118;
vmem[7667] = 8'd101;
vmem[7668] = 8'd108;
vmem[7669] = 8'd105;
vmem[7670] = 8'd116;
vmem[7671] = 8'd32;
vmem[7672] = 8'd105;
vmem[7673] = 8'd100;
vmem[7674] = 8'd44;
vmem[7675] = 8'd32;
vmem[7676] = 8'd99;
vmem[7677] = 8'd111;
vmem[7678] = 8'd110;
vmem[7679] = 8'd115;
vmem[7680] = 8'd101;
vmem[7681] = 8'd113;
vmem[7682] = 8'd117;
vmem[7683] = 8'd97;
vmem[7684] = 8'd116;
vmem[7685] = 8'd32;
vmem[7686] = 8'd111;
vmem[7687] = 8'd114;
vmem[7688] = 8'd99;
vmem[7689] = 8'd105;
vmem[7690] = 8'd46;
vmem[7691] = 8'd32;
vmem[7692] = 8'd83;
vmem[7693] = 8'd117;
vmem[7694] = 8'd115;
vmem[7695] = 8'd112;
vmem[7696] = 8'd101;
vmem[7697] = 8'd110;
vmem[7698] = 8'd100;
vmem[7699] = 8'd105;
vmem[7700] = 8'd115;
vmem[7701] = 8'd115;
vmem[7702] = 8'd101;
vmem[7703] = 8'd32;
vmem[7704] = 8'd106;
vmem[7705] = 8'd117;
vmem[7706] = 8'd115;
vmem[7707] = 8'd116;
vmem[7708] = 8'd111;
vmem[7709] = 8'd32;
vmem[7710] = 8'd109;
vmem[7711] = 8'd97;
vmem[7712] = 8'd103;
vmem[7713] = 8'd110;
vmem[7714] = 8'd97;
vmem[7715] = 8'd44;
vmem[7716] = 8'd32;
vmem[7717] = 8'd102;
vmem[7718] = 8'd101;
vmem[7719] = 8'd114;
vmem[7720] = 8'd109;
vmem[7721] = 8'd101;
vmem[7722] = 8'd110;
vmem[7723] = 8'd116;
vmem[7724] = 8'd117;
vmem[7725] = 8'd109;
vmem[7726] = 8'd32;
vmem[7727] = 8'd110;
vmem[7728] = 8'd101;
vmem[7729] = 8'd99;
vmem[7730] = 8'd32;
vmem[7731] = 8'd99;
vmem[7732] = 8'd111;
vmem[7733] = 8'd110;
vmem[7734] = 8'd103;
vmem[7735] = 8'd117;
vmem[7736] = 8'd101;
vmem[7737] = 8'd32;
vmem[7738] = 8'd97;
vmem[7739] = 8'd44;
vmem[7740] = 8'd32;
vmem[7741] = 8'd112;
vmem[7742] = 8'd117;
vmem[7743] = 8'd108;
vmem[7744] = 8'd118;
vmem[7745] = 8'd105;
vmem[7746] = 8'd110;
vmem[7747] = 8'd97;
vmem[7748] = 8'd114;
vmem[7749] = 8'd32;
vmem[7750] = 8'd118;
vmem[7751] = 8'd105;
vmem[7752] = 8'd116;
vmem[7753] = 8'd97;
vmem[7754] = 8'd101;
vmem[7755] = 8'd32;
vmem[7756] = 8'd110;
vmem[7757] = 8'd117;
vmem[7758] = 8'd110;
vmem[7759] = 8'd99;
vmem[7760] = 8'd46;
vmem[7761] = 8'd32;
vmem[7762] = 8'd81;
vmem[7763] = 8'd117;
vmem[7764] = 8'd105;
vmem[7765] = 8'd115;
vmem[7766] = 8'd113;
vmem[7767] = 8'd117;
vmem[7768] = 8'd101;
vmem[7769] = 8'd32;
vmem[7770] = 8'd101;
vmem[7771] = 8'd108;
vmem[7772] = 8'd101;
vmem[7773] = 8'd109;
vmem[7774] = 8'd101;
vmem[7775] = 8'd110;
vmem[7776] = 8'd116;
vmem[7777] = 8'd117;
vmem[7778] = 8'd109;
vmem[7779] = 8'd32;
vmem[7780] = 8'd112;
vmem[7781] = 8'd111;
vmem[7782] = 8'd115;
vmem[7783] = 8'd117;
vmem[7784] = 8'd101;
vmem[7785] = 8'd114;
vmem[7786] = 8'd101;
vmem[7787] = 8'd32;
vmem[7788] = 8'd108;
vmem[7789] = 8'd105;
vmem[7790] = 8'd103;
vmem[7791] = 8'd117;
vmem[7792] = 8'd108;
vmem[7793] = 8'd97;
vmem[7794] = 8'd32;
vmem[7795] = 8'd118;
vmem[7796] = 8'd101;
vmem[7797] = 8'd108;
vmem[7798] = 8'd32;
vmem[7799] = 8'd116;
vmem[7800] = 8'd114;
vmem[7801] = 8'd105;
vmem[7802] = 8'd115;
vmem[7803] = 8'd116;
vmem[7804] = 8'd105;
vmem[7805] = 8'd113;
vmem[7806] = 8'd117;
vmem[7807] = 8'd101;
vmem[7808] = 8'd46;
vmem[7809] = 8'd32;
vmem[7810] = 8'd83;
vmem[7811] = 8'd117;
vmem[7812] = 8'd115;
vmem[7813] = 8'd112;
vmem[7814] = 8'd101;
vmem[7815] = 8'd110;
vmem[7816] = 8'd100;
vmem[7817] = 8'd105;
vmem[7818] = 8'd115;
vmem[7819] = 8'd115;
vmem[7820] = 8'd101;
vmem[7821] = 8'd32;
vmem[7822] = 8'd98;
vmem[7823] = 8'd105;
vmem[7824] = 8'd98;
vmem[7825] = 8'd101;
vmem[7826] = 8'd110;
vmem[7827] = 8'd100;
vmem[7828] = 8'd117;
vmem[7829] = 8'd109;
vmem[7830] = 8'd32;
vmem[7831] = 8'd112;
vmem[7832] = 8'd111;
vmem[7833] = 8'd114;
vmem[7834] = 8'd116;
vmem[7835] = 8'd116;
vmem[7836] = 8'd105;
vmem[7837] = 8'd116;
vmem[7838] = 8'd111;
vmem[7839] = 8'd114;
vmem[7840] = 8'd32;
vmem[7841] = 8'd106;
vmem[7842] = 8'd117;
vmem[7843] = 8'd115;
vmem[7844] = 8'd116;
vmem[7845] = 8'd111;
vmem[7846] = 8'd32;
vmem[7847] = 8'd101;
vmem[7848] = 8'd116;
vmem[7849] = 8'd32;
vmem[7850] = 8'd116;
vmem[7851] = 8'd105;
vmem[7852] = 8'd110;
vmem[7853] = 8'd99;
vmem[7854] = 8'd105;
vmem[7855] = 8'd100;
vmem[7856] = 8'd117;
vmem[7857] = 8'd110;
vmem[7858] = 8'd116;
vmem[7859] = 8'd46;
vmem[7860] = 8'd32;
vmem[7861] = 8'd68;
vmem[7862] = 8'd111;
vmem[7863] = 8'd110;
vmem[7864] = 8'd101;
vmem[7865] = 8'd99;
vmem[7866] = 8'd32;
vmem[7867] = 8'd101;
vmem[7868] = 8'd103;
vmem[7869] = 8'd101;
vmem[7870] = 8'd116;
vmem[7871] = 8'd32;
vmem[7872] = 8'd105;
vmem[7873] = 8'd109;
vmem[7874] = 8'd112;
vmem[7875] = 8'd101;
vmem[7876] = 8'd114;
vmem[7877] = 8'd100;
vmem[7878] = 8'd105;
vmem[7879] = 8'd101;
vmem[7880] = 8'd116;
vmem[7881] = 8'd32;
vmem[7882] = 8'd100;
vmem[7883] = 8'd105;
vmem[7884] = 8'd97;
vmem[7885] = 8'd109;
vmem[7886] = 8'd44;
vmem[7887] = 8'd32;
vmem[7888] = 8'd97;
vmem[7889] = 8'd32;
vmem[7890] = 8'd102;
vmem[7891] = 8'd114;
vmem[7892] = 8'd105;
vmem[7893] = 8'd110;
vmem[7894] = 8'd103;
vmem[7895] = 8'd105;
vmem[7896] = 8'd108;
vmem[7897] = 8'd108;
vmem[7898] = 8'd97;
vmem[7899] = 8'd32;
vmem[7900] = 8'd110;
vmem[7901] = 8'd105;
vmem[7902] = 8'd115;
vmem[7903] = 8'd105;
vmem[7904] = 8'd46;
vmem[7905] = 8'd32;
vmem[7906] = 8'd65;
vmem[7907] = 8'd108;
vmem[7908] = 8'd105;
vmem[7909] = 8'd113;
vmem[7910] = 8'd117;
vmem[7911] = 8'd97;
vmem[7912] = 8'd109;
vmem[7913] = 8'd32;
vmem[7914] = 8'd101;
vmem[7915] = 8'd114;
vmem[7916] = 8'd97;
vmem[7917] = 8'd116;
vmem[7918] = 8'd32;
vmem[7919] = 8'd118;
vmem[7920] = 8'd111;
vmem[7921] = 8'd108;
vmem[7922] = 8'd117;
vmem[7923] = 8'd116;
vmem[7924] = 8'd112;
vmem[7925] = 8'd97;
vmem[7926] = 8'd116;
vmem[7927] = 8'd46;
vmem[7928] = 8'd32;
vmem[7929] = 8'd67;
vmem[7930] = 8'd117;
vmem[7931] = 8'd114;
vmem[7932] = 8'd97;
vmem[7933] = 8'd98;
vmem[7934] = 8'd105;
vmem[7935] = 8'd116;
vmem[7936] = 8'd117;
vmem[7937] = 8'd114;
vmem[7938] = 8'd32;
vmem[7939] = 8'd105;
vmem[7940] = 8'd109;
vmem[7941] = 8'd112;
vmem[7942] = 8'd101;
vmem[7943] = 8'd114;
vmem[7944] = 8'd100;
vmem[7945] = 8'd105;
vmem[7946] = 8'd101;
vmem[7947] = 8'd116;
vmem[7948] = 8'd32;
vmem[7949] = 8'd101;
vmem[7950] = 8'd115;
vmem[7951] = 8'd116;
vmem[7952] = 8'd32;
vmem[7953] = 8'd118;
vmem[7954] = 8'd101;
vmem[7955] = 8'd108;
vmem[7956] = 8'd32;
vmem[7957] = 8'd109;
vmem[7958] = 8'd105;
vmem[7959] = 8'd32;
vmem[7960] = 8'd112;
vmem[7961] = 8'd104;
vmem[7962] = 8'd97;
vmem[7963] = 8'd114;
vmem[7964] = 8'd101;
vmem[7965] = 8'd116;
vmem[7966] = 8'd114;
vmem[7967] = 8'd97;
vmem[7968] = 8'd32;
vmem[7969] = 8'd108;
vmem[7970] = 8'd97;
vmem[7971] = 8'd111;
vmem[7972] = 8'd114;
vmem[7973] = 8'd101;
vmem[7974] = 8'd101;
vmem[7975] = 8'd116;
vmem[7976] = 8'd46;
vmem[7977] = 8'd32;
vmem[7978] = 8'd80;
vmem[7979] = 8'd101;
vmem[7980] = 8'd108;
vmem[7981] = 8'd108;
vmem[7982] = 8'd101;
vmem[7983] = 8'd110;
vmem[7984] = 8'd116;
vmem[7985] = 8'd101;
vmem[7986] = 8'd115;
vmem[7987] = 8'd113;
vmem[7988] = 8'd117;
vmem[7989] = 8'd101;
vmem[7990] = 8'd32;
vmem[7991] = 8'd100;
vmem[7992] = 8'd105;
vmem[7993] = 8'd99;
vmem[7994] = 8'd116;
vmem[7995] = 8'd117;
vmem[7996] = 8'd109;
vmem[7997] = 8'd32;
vmem[7998] = 8'd97;
vmem[7999] = 8'd117;
vmem[8000] = 8'd99;
vmem[8001] = 8'd116;
vmem[8002] = 8'd111;
vmem[8003] = 8'd114;
vmem[8004] = 8'd32;
vmem[8005] = 8'd108;
vmem[8006] = 8'd101;
vmem[8007] = 8'd99;
vmem[8008] = 8'd116;
vmem[8009] = 8'd117;
vmem[8010] = 8'd115;
vmem[8011] = 8'd44;
vmem[8012] = 8'd32;
vmem[8013] = 8'd101;
vmem[8014] = 8'd108;
vmem[8015] = 8'd101;
vmem[8016] = 8'd109;
vmem[8017] = 8'd101;
vmem[8018] = 8'd110;
vmem[8019] = 8'd116;
vmem[8020] = 8'd117;
vmem[8021] = 8'd109;
vmem[8022] = 8'd32;
vmem[8023] = 8'd112;
vmem[8024] = 8'd111;
vmem[8025] = 8'd114;
vmem[8026] = 8'd116;
vmem[8027] = 8'd116;
vmem[8028] = 8'd105;
vmem[8029] = 8'd116;
vmem[8030] = 8'd111;
vmem[8031] = 8'd114;
vmem[8032] = 8'd32;
vmem[8033] = 8'd100;
vmem[8034] = 8'd117;
vmem[8035] = 8'd105;
vmem[8036] = 8'd32;
vmem[8037] = 8'd102;
vmem[8038] = 8'd97;
vmem[8039] = 8'd117;
vmem[8040] = 8'd99;
vmem[8041] = 8'd105;
vmem[8042] = 8'd98;
vmem[8043] = 8'd117;
vmem[8044] = 8'd115;
vmem[8045] = 8'd32;
vmem[8046] = 8'd118;
vmem[8047] = 8'd97;
vmem[8048] = 8'd114;
vmem[8049] = 8'd105;
vmem[8050] = 8'd117;
vmem[8051] = 8'd115;
vmem[8052] = 8'd46;
vmem[8053] = 8'd32;
vmem[8054] = 8'd80;
vmem[8055] = 8'd101;
vmem[8056] = 8'd108;
vmem[8057] = 8'd108;
vmem[8058] = 8'd101;
vmem[8059] = 8'd110;
vmem[8060] = 8'd116;
vmem[8061] = 8'd101;
vmem[8062] = 8'd115;
vmem[8063] = 8'd113;
vmem[8064] = 8'd117;
vmem[8065] = 8'd101;
vmem[8066] = 8'd32;
vmem[8067] = 8'd116;
vmem[8068] = 8'd101;
vmem[8069] = 8'd109;
vmem[8070] = 8'd112;
vmem[8071] = 8'd111;
vmem[8072] = 8'd114;
vmem[8073] = 8'd32;
vmem[8074] = 8'd108;
vmem[8075] = 8'd97;
vmem[8076] = 8'd99;
vmem[8077] = 8'd105;
vmem[8078] = 8'd110;
vmem[8079] = 8'd105;
vmem[8080] = 8'd97;
vmem[8081] = 8'd32;
vmem[8082] = 8'd108;
vmem[8083] = 8'd101;
vmem[8084] = 8'd99;
vmem[8085] = 8'd116;
vmem[8086] = 8'd117;
vmem[8087] = 8'd115;
vmem[8088] = 8'd32;
vmem[8089] = 8'd101;
vmem[8090] = 8'd116;
vmem[8091] = 8'd32;
vmem[8092] = 8'd118;
vmem[8093] = 8'd97;
vmem[8094] = 8'd114;
vmem[8095] = 8'd105;
vmem[8096] = 8'd117;
vmem[8097] = 8'd115;
vmem[8098] = 8'd46;
vmem[8099] = 8'd32;
vmem[8100] = 8'd69;
vmem[8101] = 8'd116;
vmem[8102] = 8'd105;
vmem[8103] = 8'd97;
vmem[8104] = 8'd109;
vmem[8105] = 8'd32;
vmem[8106] = 8'd97;
vmem[8107] = 8'd32;
vmem[8108] = 8'd100;
vmem[8109] = 8'd105;
vmem[8110] = 8'd97;
vmem[8111] = 8'd109;
vmem[8112] = 8'd32;
vmem[8113] = 8'd118;
vmem[8114] = 8'd111;
vmem[8115] = 8'd108;
vmem[8116] = 8'd117;
vmem[8117] = 8'd116;
vmem[8118] = 8'd112;
vmem[8119] = 8'd97;
vmem[8120] = 8'd116;
vmem[8121] = 8'd44;
vmem[8122] = 8'd32;
vmem[8123] = 8'd112;
vmem[8124] = 8'd101;
vmem[8125] = 8'd108;
vmem[8126] = 8'd108;
vmem[8127] = 8'd101;
vmem[8128] = 8'd110;
vmem[8129] = 8'd116;
vmem[8130] = 8'd101;
vmem[8131] = 8'd115;
vmem[8132] = 8'd113;
vmem[8133] = 8'd117;
vmem[8134] = 8'd101;
vmem[8135] = 8'd32;
vmem[8136] = 8'd108;
vmem[8137] = 8'd111;
vmem[8138] = 8'd114;
vmem[8139] = 8'd101;
vmem[8140] = 8'd109;
vmem[8141] = 8'd32;
vmem[8142] = 8'd97;
vmem[8143] = 8'd99;
vmem[8144] = 8'd44;
vmem[8145] = 8'd32;
vmem[8146] = 8'd97;
vmem[8147] = 8'd108;
vmem[8148] = 8'd105;
vmem[8149] = 8'd113;
vmem[8150] = 8'd117;
vmem[8151] = 8'd97;
vmem[8152] = 8'd109;
vmem[8153] = 8'd32;
vmem[8154] = 8'd101;
vmem[8155] = 8'd108;
vmem[8156] = 8'd105;
vmem[8157] = 8'd116;
vmem[8158] = 8'd46;
vmem[8159] = 8'd32;
vmem[8160] = 8'd68;
vmem[8161] = 8'd117;
vmem[8162] = 8'd105;
vmem[8163] = 8'd115;
vmem[8164] = 8'd32;
vmem[8165] = 8'd114;
vmem[8166] = 8'd117;
vmem[8167] = 8'd116;
vmem[8168] = 8'd114;
vmem[8169] = 8'd117;
vmem[8170] = 8'd109;
vmem[8171] = 8'd44;
vmem[8172] = 8'd32;
vmem[8173] = 8'd110;
vmem[8174] = 8'd101;
vmem[8175] = 8'd113;
vmem[8176] = 8'd117;
vmem[8177] = 8'd101;
vmem[8178] = 8'd32;
vmem[8179] = 8'd97;
vmem[8180] = 8'd32;
vmem[8181] = 8'd111;
vmem[8182] = 8'd114;
vmem[8183] = 8'd110;
vmem[8184] = 8'd97;
vmem[8185] = 8'd114;
vmem[8186] = 8'd101;
vmem[8187] = 8'd32;
vmem[8188] = 8'd108;
vmem[8189] = 8'd117;
vmem[8190] = 8'd99;
vmem[8191] = 8'd116;
vmem[8192] = 8'd117;
vmem[8193] = 8'd115;
vmem[8194] = 8'd44;
vmem[8195] = 8'd32;
vmem[8196] = 8'd101;
vmem[8197] = 8'd110;
vmem[8198] = 8'd105;
vmem[8199] = 8'd109;
vmem[8200] = 8'd32;
vmem[8201] = 8'd116;
vmem[8202] = 8'd117;
vmem[8203] = 8'd114;
vmem[8204] = 8'd112;
vmem[8205] = 8'd105;
vmem[8206] = 8'd115;
vmem[8207] = 8'd32;
vmem[8208] = 8'd116;
vmem[8209] = 8'd114;
vmem[8210] = 8'd105;
vmem[8211] = 8'd115;
vmem[8212] = 8'd116;
vmem[8213] = 8'd105;
vmem[8214] = 8'd113;
vmem[8215] = 8'd117;
vmem[8216] = 8'd101;
vmem[8217] = 8'd32;
vmem[8218] = 8'd113;
vmem[8219] = 8'd117;
vmem[8220] = 8'd97;
vmem[8221] = 8'd109;
vmem[8222] = 8'd44;
vmem[8223] = 8'd32;
vmem[8224] = 8'd118;
vmem[8225] = 8'd105;
vmem[8226] = 8'd116;
vmem[8227] = 8'd97;
vmem[8228] = 8'd101;
vmem[8229] = 8'd32;
vmem[8230] = 8'd102;
vmem[8231] = 8'd101;
vmem[8232] = 8'd117;
vmem[8233] = 8'd103;
vmem[8234] = 8'd105;
vmem[8235] = 8'd97;
vmem[8236] = 8'd116;
vmem[8237] = 8'd32;
vmem[8238] = 8'd101;
vmem[8239] = 8'd114;
vmem[8240] = 8'd97;
vmem[8241] = 8'd116;
vmem[8242] = 8'd32;
vmem[8243] = 8'd102;
vmem[8244] = 8'd101;
vmem[8245] = 8'd108;
vmem[8246] = 8'd105;
vmem[8247] = 8'd115;
vmem[8248] = 8'd32;
vmem[8249] = 8'd97;
vmem[8250] = 8'd99;
vmem[8251] = 8'd32;
vmem[8252] = 8'd110;
vmem[8253] = 8'd101;
vmem[8254] = 8'd113;
vmem[8255] = 8'd117;
vmem[8256] = 8'd101;
vmem[8257] = 8'd46;
vmem[8258] = 8'd32;
vmem[8259] = 8'd68;
vmem[8260] = 8'd117;
vmem[8261] = 8'd105;
vmem[8262] = 8'd115;
vmem[8263] = 8'd32;
vmem[8264] = 8'd110;
vmem[8265] = 8'd101;
vmem[8266] = 8'd99;
vmem[8267] = 8'd32;
vmem[8268] = 8'd108;
vmem[8269] = 8'd97;
vmem[8270] = 8'd99;
vmem[8271] = 8'd117;
vmem[8272] = 8'd115;
vmem[8273] = 8'd32;
vmem[8274] = 8'd118;
vmem[8275] = 8'd111;
vmem[8276] = 8'd108;
vmem[8277] = 8'd117;
vmem[8278] = 8'd116;
vmem[8279] = 8'd112;
vmem[8280] = 8'd97;
vmem[8281] = 8'd116;
vmem[8282] = 8'd44;
vmem[8283] = 8'd32;
vmem[8284] = 8'd112;
vmem[8285] = 8'd111;
vmem[8286] = 8'd114;
vmem[8287] = 8'd116;
vmem[8288] = 8'd97;
vmem[8289] = 8'd32;
vmem[8290] = 8'd116;
vmem[8291] = 8'd111;
vmem[8292] = 8'd114;
vmem[8293] = 8'd116;
vmem[8294] = 8'd111;
vmem[8295] = 8'd114;
vmem[8296] = 8'd32;
vmem[8297] = 8'd97;
vmem[8298] = 8'd44;
vmem[8299] = 8'd32;
vmem[8300] = 8'd100;
vmem[8301] = 8'd97;
vmem[8302] = 8'd112;
vmem[8303] = 8'd105;
vmem[8304] = 8'd98;
vmem[8305] = 8'd117;
vmem[8306] = 8'd115;
vmem[8307] = 8'd32;
vmem[8308] = 8'd118;
vmem[8309] = 8'd101;
vmem[8310] = 8'd108;
vmem[8311] = 8'd105;
vmem[8312] = 8'd116;
vmem[8313] = 8'd46;
vmem[8314] = 8'd32;
vmem[8315] = 8'd76;
vmem[8316] = 8'd111;
vmem[8317] = 8'd114;
vmem[8318] = 8'd101;
vmem[8319] = 8'd109;
vmem[8320] = 8'd32;
vmem[8321] = 8'd105;
vmem[8322] = 8'd112;
vmem[8323] = 8'd115;
vmem[8324] = 8'd117;
vmem[8325] = 8'd109;
vmem[8326] = 8'd32;
vmem[8327] = 8'd100;
vmem[8328] = 8'd111;
vmem[8329] = 8'd108;
vmem[8330] = 8'd111;
vmem[8331] = 8'd114;
vmem[8332] = 8'd32;
vmem[8333] = 8'd115;
vmem[8334] = 8'd105;
vmem[8335] = 8'd116;
vmem[8336] = 8'd32;
vmem[8337] = 8'd97;
vmem[8338] = 8'd109;
vmem[8339] = 8'd101;
vmem[8340] = 8'd116;
vmem[8341] = 8'd44;
vmem[8342] = 8'd32;
vmem[8343] = 8'd99;
vmem[8344] = 8'd111;
vmem[8345] = 8'd110;
vmem[8346] = 8'd115;
vmem[8347] = 8'd101;
vmem[8348] = 8'd99;
vmem[8349] = 8'd116;
vmem[8350] = 8'd101;
vmem[8351] = 8'd116;
vmem[8352] = 8'd117;
vmem[8353] = 8'd114;
vmem[8354] = 8'd32;
vmem[8355] = 8'd97;
vmem[8356] = 8'd100;
vmem[8357] = 8'd105;
vmem[8358] = 8'd112;
vmem[8359] = 8'd105;
vmem[8360] = 8'd115;
vmem[8361] = 8'd99;
vmem[8362] = 8'd105;
vmem[8363] = 8'd110;
vmem[8364] = 8'd103;
vmem[8365] = 8'd32;
vmem[8366] = 8'd101;
vmem[8367] = 8'd108;
vmem[8368] = 8'd105;
vmem[8369] = 8'd116;
vmem[8370] = 8'd46;
vmem[8371] = 8'd32;
vmem[8372] = 8'd80;
vmem[8373] = 8'd101;
vmem[8374] = 8'd108;
vmem[8375] = 8'd108;
vmem[8376] = 8'd101;
vmem[8377] = 8'd110;
vmem[8378] = 8'd116;
vmem[8379] = 8'd101;
vmem[8380] = 8'd115;
vmem[8381] = 8'd113;
vmem[8382] = 8'd117;
vmem[8383] = 8'd101;
vmem[8384] = 8'd32;
vmem[8385] = 8'd115;
vmem[8386] = 8'd117;
vmem[8387] = 8'd115;
vmem[8388] = 8'd99;
vmem[8389] = 8'd105;
vmem[8390] = 8'd112;
vmem[8391] = 8'd105;
vmem[8392] = 8'd116;
vmem[8393] = 8'd32;
vmem[8394] = 8'd102;
vmem[8395] = 8'd105;
vmem[8396] = 8'd110;
vmem[8397] = 8'd105;
vmem[8398] = 8'd98;
vmem[8399] = 8'd117;
vmem[8400] = 8'd115;
vmem[8401] = 8'd32;
vmem[8402] = 8'd117;
vmem[8403] = 8'd108;
vmem[8404] = 8'd116;
vmem[8405] = 8'd114;
vmem[8406] = 8'd105;
vmem[8407] = 8'd99;
vmem[8408] = 8'd101;
vmem[8409] = 8'd115;
vmem[8410] = 8'd46;
vmem[8411] = 8'd32;
vmem[8412] = 8'd86;
vmem[8413] = 8'd105;
vmem[8414] = 8'd118;
vmem[8415] = 8'd97;
vmem[8416] = 8'd109;
vmem[8417] = 8'd117;
vmem[8418] = 8'd115;
vmem[8419] = 8'd32;
vmem[8420] = 8'd99;
vmem[8421] = 8'd111;
vmem[8422] = 8'd109;
vmem[8423] = 8'd109;
vmem[8424] = 8'd111;
vmem[8425] = 8'd100;
vmem[8426] = 8'd111;
vmem[8427] = 8'd32;
vmem[8428] = 8'd109;
vmem[8429] = 8'd105;
vmem[8430] = 8'd32;
vmem[8431] = 8'd102;
vmem[8432] = 8'd101;
vmem[8433] = 8'd108;
vmem[8434] = 8'd105;
vmem[8435] = 8'd115;
vmem[8436] = 8'd46;
vmem[8437] = 8'd32;
vmem[8438] = 8'd83;
vmem[8439] = 8'd101;
vmem[8440] = 8'd100;
vmem[8441] = 8'd32;
vmem[8442] = 8'd110;
vmem[8443] = 8'd111;
vmem[8444] = 8'd110;
vmem[8445] = 8'd32;
vmem[8446] = 8'd117;
vmem[8447] = 8'd108;
vmem[8448] = 8'd116;
vmem[8449] = 8'd114;
vmem[8450] = 8'd105;
vmem[8451] = 8'd99;
vmem[8452] = 8'd101;
vmem[8453] = 8'd115;
vmem[8454] = 8'd32;
vmem[8455] = 8'd109;
vmem[8456] = 8'd105;
vmem[8457] = 8'd46;
vmem[8458] = 8'd32;
vmem[8459] = 8'd68;
vmem[8460] = 8'd117;
vmem[8461] = 8'd105;
vmem[8462] = 8'd115;
vmem[8463] = 8'd32;
vmem[8464] = 8'd114;
vmem[8465] = 8'd104;
vmem[8466] = 8'd111;
vmem[8467] = 8'd110;
vmem[8468] = 8'd99;
vmem[8469] = 8'd117;
vmem[8470] = 8'd115;
vmem[8471] = 8'd44;
vmem[8472] = 8'd32;
vmem[8473] = 8'd109;
vmem[8474] = 8'd105;
vmem[8475] = 8'd32;
vmem[8476] = 8'd105;
vmem[8477] = 8'd110;
vmem[8478] = 8'd32;
vmem[8479] = 8'd105;
vmem[8480] = 8'd97;
vmem[8481] = 8'd99;
vmem[8482] = 8'd117;
vmem[8483] = 8'd108;
vmem[8484] = 8'd105;
vmem[8485] = 8'd115;
vmem[8486] = 8'd32;
vmem[8487] = 8'd109;
vmem[8488] = 8'd97;
vmem[8489] = 8'd116;
vmem[8490] = 8'd116;
vmem[8491] = 8'd105;
vmem[8492] = 8'd115;
vmem[8493] = 8'd44;
vmem[8494] = 8'd32;
vmem[8495] = 8'd101;
vmem[8496] = 8'd120;
vmem[8497] = 8'd32;
vmem[8498] = 8'd100;
vmem[8499] = 8'd117;
vmem[8500] = 8'd105;
vmem[8501] = 8'd32;
vmem[8502] = 8'd118;
vmem[8503] = 8'd101;
vmem[8504] = 8'd110;
vmem[8505] = 8'd101;
vmem[8506] = 8'd110;
vmem[8507] = 8'd97;
vmem[8508] = 8'd116;
vmem[8509] = 8'd105;
vmem[8510] = 8'd115;
vmem[8511] = 8'd32;
vmem[8512] = 8'd111;
vmem[8513] = 8'd100;
vmem[8514] = 8'd105;
vmem[8515] = 8'd111;
vmem[8516] = 8'd44;
vmem[8517] = 8'd32;
vmem[8518] = 8'd105;
vmem[8519] = 8'd100;
vmem[8520] = 8'd32;
vmem[8521] = 8'd99;
vmem[8522] = 8'd117;
vmem[8523] = 8'd114;
vmem[8524] = 8'd115;
vmem[8525] = 8'd117;
vmem[8526] = 8'd115;
vmem[8527] = 8'd32;
vmem[8528] = 8'd108;
vmem[8529] = 8'd101;
vmem[8530] = 8'd111;
vmem[8531] = 8'd32;
vmem[8532] = 8'd116;
vmem[8533] = 8'd117;
vmem[8534] = 8'd114;
vmem[8535] = 8'd112;
vmem[8536] = 8'd105;
vmem[8537] = 8'd115;
vmem[8538] = 8'd32;
vmem[8539] = 8'd99;
vmem[8540] = 8'd111;
vmem[8541] = 8'd110;
vmem[8542] = 8'd103;
vmem[8543] = 8'd117;
vmem[8544] = 8'd101;
vmem[8545] = 8'd32;
vmem[8546] = 8'd101;
vmem[8547] = 8'd114;
vmem[8548] = 8'd111;
vmem[8549] = 8'd115;
vmem[8550] = 8'd46;
vmem[8551] = 8'd32;
vmem[8552] = 8'd86;
vmem[8553] = 8'd105;
vmem[8554] = 8'd118;
vmem[8555] = 8'd97;
vmem[8556] = 8'd109;
vmem[8557] = 8'd117;
vmem[8558] = 8'd115;
vmem[8559] = 8'd32;
vmem[8560] = 8'd101;
vmem[8561] = 8'd103;
vmem[8562] = 8'd101;
vmem[8563] = 8'd116;
vmem[8564] = 8'd32;
vmem[8565] = 8'd109;
vmem[8566] = 8'd97;
vmem[8567] = 8'd115;
vmem[8568] = 8'd115;
vmem[8569] = 8'd97;
vmem[8570] = 8'd32;
vmem[8571] = 8'd110;
vmem[8572] = 8'd101;
vmem[8573] = 8'd99;
vmem[8574] = 8'd32;
vmem[8575] = 8'd108;
vmem[8576] = 8'd101;
vmem[8577] = 8'd99;
vmem[8578] = 8'd116;
vmem[8579] = 8'd117;
vmem[8580] = 8'd115;
vmem[8581] = 8'd32;
vmem[8582] = 8'd112;
vmem[8583] = 8'd101;
vmem[8584] = 8'd108;
vmem[8585] = 8'd108;
vmem[8586] = 8'd101;
vmem[8587] = 8'd110;
vmem[8588] = 8'd116;
vmem[8589] = 8'd101;
vmem[8590] = 8'd115;
vmem[8591] = 8'd113;
vmem[8592] = 8'd117;
vmem[8593] = 8'd101;
vmem[8594] = 8'd32;
vmem[8595] = 8'd117;
vmem[8596] = 8'd108;
vmem[8597] = 8'd116;
vmem[8598] = 8'd114;
vmem[8599] = 8'd105;
vmem[8600] = 8'd99;
vmem[8601] = 8'd105;
vmem[8602] = 8'd101;
vmem[8603] = 8'd115;
vmem[8604] = 8'd46;
vmem[8605] = 8'd32;
vmem[8606] = 8'd77;
vmem[8607] = 8'd97;
vmem[8608] = 8'd101;
vmem[8609] = 8'd99;
vmem[8610] = 8'd101;
vmem[8611] = 8'd110;
vmem[8612] = 8'd97;
vmem[8613] = 8'd115;
vmem[8614] = 8'd32;
vmem[8615] = 8'd97;
vmem[8616] = 8'd108;
vmem[8617] = 8'd105;
vmem[8618] = 8'd113;
vmem[8619] = 8'd117;
vmem[8620] = 8'd97;
vmem[8621] = 8'd109;
vmem[8622] = 8'd32;
vmem[8623] = 8'd115;
vmem[8624] = 8'd97;
vmem[8625] = 8'd112;
vmem[8626] = 8'd105;
vmem[8627] = 8'd101;
vmem[8628] = 8'd110;
vmem[8629] = 8'd32;
vmem[8630] = 8'd118;
vmem[8631] = 8'd101;
vmem[8632] = 8'd108;
vmem[8633] = 8'd32;
vmem[8634] = 8'd112;
vmem[8635] = 8'd108;
vmem[8636] = 8'd97;
vmem[8637] = 8'd99;
vmem[8638] = 8'd101;
vmem[8639] = 8'd114;
vmem[8640] = 8'd97;
vmem[8641] = 8'd116;
vmem[8642] = 8'd32;
vmem[8643] = 8'd97;
vmem[8644] = 8'd117;
vmem[8645] = 8'd99;
vmem[8646] = 8'd116;
vmem[8647] = 8'd111;
vmem[8648] = 8'd114;
vmem[8649] = 8'd46;
vmem[8650] = 8'd32;
vmem[8651] = 8'd85;
vmem[8652] = 8'd116;
vmem[8653] = 8'd32;
vmem[8654] = 8'd109;
vmem[8655] = 8'd111;
vmem[8656] = 8'd108;
vmem[8657] = 8'd108;
vmem[8658] = 8'd105;
vmem[8659] = 8'd115;
vmem[8660] = 8'd32;
vmem[8661] = 8'd97;
vmem[8662] = 8'd99;
vmem[8663] = 8'd32;
vmem[8664] = 8'd102;
vmem[8665] = 8'd101;
vmem[8666] = 8'd108;
vmem[8667] = 8'd105;
vmem[8668] = 8'd115;
vmem[8669] = 8'd32;
vmem[8670] = 8'd110;
vmem[8671] = 8'd101;
vmem[8672] = 8'd99;
vmem[8673] = 8'd32;
vmem[8674] = 8'd118;
vmem[8675] = 8'd101;
vmem[8676] = 8'd110;
vmem[8677] = 8'd101;
vmem[8678] = 8'd110;
vmem[8679] = 8'd97;
vmem[8680] = 8'd116;
vmem[8681] = 8'd105;
vmem[8682] = 8'd115;
vmem[8683] = 8'd46;
vmem[8684] = 8'd32;
vmem[8685] = 8'd68;
vmem[8686] = 8'd117;
vmem[8687] = 8'd105;
vmem[8688] = 8'd115;
vmem[8689] = 8'd32;
vmem[8690] = 8'd115;
vmem[8691] = 8'd101;
vmem[8692] = 8'd100;
vmem[8693] = 8'd32;
vmem[8694] = 8'd109;
vmem[8695] = 8'd97;
vmem[8696] = 8'd103;
vmem[8697] = 8'd110;
vmem[8698] = 8'd97;
vmem[8699] = 8'd32;
vmem[8700] = 8'd118;
vmem[8701] = 8'd105;
vmem[8702] = 8'd118;
vmem[8703] = 8'd101;
vmem[8704] = 8'd114;
vmem[8705] = 8'd114;
vmem[8706] = 8'd97;
vmem[8707] = 8'd44;
vmem[8708] = 8'd32;
vmem[8709] = 8'd112;
vmem[8710] = 8'd108;
vmem[8711] = 8'd97;
vmem[8712] = 8'd99;
vmem[8713] = 8'd101;
vmem[8714] = 8'd114;
vmem[8715] = 8'd97;
vmem[8716] = 8'd116;
vmem[8717] = 8'd32;
vmem[8718] = 8'd101;
vmem[8719] = 8'd108;
vmem[8720] = 8'd105;
vmem[8721] = 8'd116;
vmem[8722] = 8'd32;
vmem[8723] = 8'd110;
vmem[8724] = 8'd101;
vmem[8725] = 8'd99;
vmem[8726] = 8'd44;
vmem[8727] = 8'd32;
vmem[8728] = 8'd100;
vmem[8729] = 8'd105;
vmem[8730] = 8'd99;
vmem[8731] = 8'd116;
vmem[8732] = 8'd117;
vmem[8733] = 8'd109;
vmem[8734] = 8'd32;
vmem[8735] = 8'd115;
vmem[8736] = 8'd97;
vmem[8737] = 8'd112;
vmem[8738] = 8'd105;
vmem[8739] = 8'd101;
vmem[8740] = 8'd110;
vmem[8741] = 8'd46;
vmem[8742] = 8'd32;
vmem[8743] = 8'd80;
vmem[8744] = 8'd114;
vmem[8745] = 8'd111;
vmem[8746] = 8'd105;
vmem[8747] = 8'd110;
vmem[8748] = 8'd32;
vmem[8749] = 8'd118;
vmem[8750] = 8'd101;
vmem[8751] = 8'd110;
vmem[8752] = 8'd101;
vmem[8753] = 8'd110;
vmem[8754] = 8'd97;
vmem[8755] = 8'd116;
vmem[8756] = 8'd105;
vmem[8757] = 8'd115;
vmem[8758] = 8'd32;
vmem[8759] = 8'd101;
vmem[8760] = 8'd103;
vmem[8761] = 8'd101;
vmem[8762] = 8'd115;
vmem[8763] = 8'd116;
vmem[8764] = 8'd97;
vmem[8765] = 8'd115;
vmem[8766] = 8'd32;
vmem[8767] = 8'd108;
vmem[8768] = 8'd105;
vmem[8769] = 8'd98;
vmem[8770] = 8'd101;
vmem[8771] = 8'd114;
vmem[8772] = 8'd111;
vmem[8773] = 8'd32;
vmem[8774] = 8'd97;
vmem[8775] = 8'd116;
vmem[8776] = 8'd32;
vmem[8777] = 8'd103;
vmem[8778] = 8'd114;
vmem[8779] = 8'd97;
vmem[8780] = 8'd118;
vmem[8781] = 8'd105;
vmem[8782] = 8'd100;
vmem[8783] = 8'd97;
vmem[8784] = 8'd46;
vmem[8785] = 8'd32;
vmem[8786] = 8'd77;
vmem[8787] = 8'd97;
vmem[8788] = 8'd101;
vmem[8789] = 8'd99;
vmem[8790] = 8'd101;
vmem[8791] = 8'd110;
vmem[8792] = 8'd97;
vmem[8793] = 8'd115;
vmem[8794] = 8'd32;
vmem[8795] = 8'd97;
vmem[8796] = 8'd108;
vmem[8797] = 8'd105;
vmem[8798] = 8'd113;
vmem[8799] = 8'd117;
vmem[8800] = 8'd101;
vmem[8801] = 8'd116;
vmem[8802] = 8'd32;
vmem[8803] = 8'd116;
vmem[8804] = 8'd117;
vmem[8805] = 8'd114;
vmem[8806] = 8'd112;
vmem[8807] = 8'd105;
vmem[8808] = 8'd115;
vmem[8809] = 8'd32;
vmem[8810] = 8'd105;
vmem[8811] = 8'd110;
vmem[8812] = 8'd32;
vmem[8813] = 8'd101;
vmem[8814] = 8'd115;
vmem[8815] = 8'd116;
vmem[8816] = 8'd32;
vmem[8817] = 8'd115;
vmem[8818] = 8'd111;
vmem[8819] = 8'd100;
vmem[8820] = 8'd97;
vmem[8821] = 8'd108;
vmem[8822] = 8'd101;
vmem[8823] = 8'd115;
vmem[8824] = 8'd44;
vmem[8825] = 8'd32;
vmem[8826] = 8'd105;
vmem[8827] = 8'd100;
vmem[8828] = 8'd32;
vmem[8829] = 8'd115;
vmem[8830] = 8'd97;
vmem[8831] = 8'd103;
vmem[8832] = 8'd105;
vmem[8833] = 8'd116;
vmem[8834] = 8'd116;
vmem[8835] = 8'd105;
vmem[8836] = 8'd115;
vmem[8837] = 8'd32;
vmem[8838] = 8'd116;
vmem[8839] = 8'd111;
vmem[8840] = 8'd114;
vmem[8841] = 8'd116;
vmem[8842] = 8'd111;
vmem[8843] = 8'd114;
vmem[8844] = 8'd32;
vmem[8845] = 8'd112;
vmem[8846] = 8'd111;
vmem[8847] = 8'd115;
vmem[8848] = 8'd117;
vmem[8849] = 8'd101;
vmem[8850] = 8'd114;
vmem[8851] = 8'd101;
vmem[8852] = 8'd46;
vmem[8853] = 8'd32;
vmem[8854] = 8'd77;
vmem[8855] = 8'd111;
vmem[8856] = 8'd114;
vmem[8857] = 8'd98;
vmem[8858] = 8'd105;
vmem[8859] = 8'd32;
vmem[8860] = 8'd97;
vmem[8861] = 8'd116;
vmem[8862] = 8'd32;
vmem[8863] = 8'd117;
vmem[8864] = 8'd114;
vmem[8865] = 8'd110;
vmem[8866] = 8'd97;
vmem[8867] = 8'd32;
vmem[8868] = 8'd116;
vmem[8869] = 8'd105;
vmem[8870] = 8'd110;
vmem[8871] = 8'd99;
vmem[8872] = 8'd105;
vmem[8873] = 8'd100;
vmem[8874] = 8'd117;
vmem[8875] = 8'd110;
vmem[8876] = 8'd116;
vmem[8877] = 8'd44;
vmem[8878] = 8'd32;
vmem[8879] = 8'd99;
vmem[8880] = 8'd111;
vmem[8881] = 8'd110;
vmem[8882] = 8'd115;
vmem[8883] = 8'd101;
vmem[8884] = 8'd99;
vmem[8885] = 8'd116;
vmem[8886] = 8'd101;
vmem[8887] = 8'd116;
vmem[8888] = 8'd117;
vmem[8889] = 8'd114;
vmem[8890] = 8'd32;
vmem[8891] = 8'd97;
vmem[8892] = 8'd114;
vmem[8893] = 8'd99;
vmem[8894] = 8'd117;
vmem[8895] = 8'd32;
vmem[8896] = 8'd97;
vmem[8897] = 8'd99;
vmem[8898] = 8'd44;
vmem[8899] = 8'd32;
vmem[8900] = 8'd103;
vmem[8901] = 8'd114;
vmem[8902] = 8'd97;
vmem[8903] = 8'd118;
vmem[8904] = 8'd105;
vmem[8905] = 8'd100;
vmem[8906] = 8'd97;
vmem[8907] = 8'd32;
vmem[8908] = 8'd113;
vmem[8909] = 8'd117;
vmem[8910] = 8'd97;
vmem[8911] = 8'd109;
vmem[8912] = 8'd46;
vmem[8913] = 8'd32;
vmem[8914] = 8'd77;
vmem[8915] = 8'd97;
vmem[8916] = 8'd101;
vmem[8917] = 8'd99;
vmem[8918] = 8'd101;
vmem[8919] = 8'd110;
vmem[8920] = 8'd97;
vmem[8921] = 8'd115;
vmem[8922] = 8'd32;
vmem[8923] = 8'd102;
vmem[8924] = 8'd97;
vmem[8925] = 8'd99;
vmem[8926] = 8'd105;
vmem[8927] = 8'd108;
vmem[8928] = 8'd105;
vmem[8929] = 8'd115;
vmem[8930] = 8'd105;
vmem[8931] = 8'd115;
vmem[8932] = 8'd32;
vmem[8933] = 8'd115;
vmem[8934] = 8'd97;
vmem[8935] = 8'd103;
vmem[8936] = 8'd105;
vmem[8937] = 8'd116;
vmem[8938] = 8'd116;
vmem[8939] = 8'd105;
vmem[8940] = 8'd115;
vmem[8941] = 8'd32;
vmem[8942] = 8'd108;
vmem[8943] = 8'd101;
vmem[8944] = 8'd111;
vmem[8945] = 8'd32;
vmem[8946] = 8'd105;
vmem[8947] = 8'd100;
vmem[8948] = 8'd32;
vmem[8949] = 8'd98;
vmem[8950] = 8'd108;
vmem[8951] = 8'd97;
vmem[8952] = 8'd110;
vmem[8953] = 8'd100;
vmem[8954] = 8'd105;
vmem[8955] = 8'd116;
vmem[8956] = 8'd46;
vmem[8957] = 8'd32;
vmem[8958] = 8'd77;
vmem[8959] = 8'd97;
vmem[8960] = 8'd101;
vmem[8961] = 8'd99;
vmem[8962] = 8'd101;
vmem[8963] = 8'd110;
vmem[8964] = 8'd97;
vmem[8965] = 8'd115;
vmem[8966] = 8'd32;
vmem[8967] = 8'd97;
vmem[8968] = 8'd99;
vmem[8969] = 8'd32;
vmem[8970] = 8'd109;
vmem[8971] = 8'd97;
vmem[8972] = 8'd117;
vmem[8973] = 8'd114;
vmem[8974] = 8'd105;
vmem[8975] = 8'd115;
vmem[8976] = 8'd32;
vmem[8977] = 8'd112;
vmem[8978] = 8'd111;
vmem[8979] = 8'd114;
vmem[8980] = 8'd116;
vmem[8981] = 8'd97;
vmem[8982] = 8'd32;
vmem[8983] = 8'd105;
vmem[8984] = 8'd112;
vmem[8985] = 8'd115;
vmem[8986] = 8'd117;
vmem[8987] = 8'd109;
vmem[8988] = 8'd32;
vmem[8989] = 8'd97;
vmem[8990] = 8'd99;
vmem[8991] = 8'd99;
vmem[8992] = 8'd117;
vmem[8993] = 8'd109;
vmem[8994] = 8'd115;
vmem[8995] = 8'd97;
vmem[8996] = 8'd110;
vmem[8997] = 8'd32;
vmem[8998] = 8'd101;
vmem[8999] = 8'd103;
vmem[9000] = 8'd101;
vmem[9001] = 8'd115;
vmem[9002] = 8'd116;
vmem[9003] = 8'd97;
vmem[9004] = 8'd115;
vmem[9005] = 8'd32;
vmem[9006] = 8'd113;
vmem[9007] = 8'd117;
vmem[9008] = 8'd105;
vmem[9009] = 8'd115;
vmem[9010] = 8'd32;
vmem[9011] = 8'd97;
vmem[9012] = 8'd116;
vmem[9013] = 8'd32;
vmem[9014] = 8'd101;
vmem[9015] = 8'd117;
vmem[9016] = 8'd46;
vmem[9017] = 8'd32;




    vmem [CH_SCREENSIZE-1] = 8'b11111111;
    vmem [CH_SCREENSIZE-3] = 8'b11111110;

end

endmodule
