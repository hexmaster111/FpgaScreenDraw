module XYDrawGenerator (
    input wire [9:0] i_hCount, i_vCount,
    output wire o_drawing,
    output wire [9:0] o_x_pixel, o_y_pixel
);
    
endmodule
